`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b/QhBR/oOzwaIZ6E7xuGaVjTIqrrrk1JJQRhGHM3PGlr0wSnnQxll/0isGyM+wjDSK9GtAlYP0OM
/PCkyb+ehw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WJYbCKycBENXWINGjywfHsrNXZknL7yjgguwmqs6OwjbxK0hf5LYRBnuDpYwQhonmgh8FspAKN7S
vBI1o5pda3s0NrnqYv/G6epYOX6UDWwAVMwCaLpfxBgAA/lPO47odG5bWak48ZfirMNoqxPrYu/X
xn6bfuLcmjfyW6TeE4M=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mW//b3sbAmqxeiGHJDCiVCvPi9GZokMwU+5dRZ6OAcIpAn4OGe3GYmtpujCuVoiFy4oJaeHTE0DN
0VSZByGuwXomWUNjVxzi6wOCqyMnHN+CyPAWgXBhdnVWIXrkwfog4y5TSHD++gZeUJPFrxmlbbwN
+DAsGPPK04f6ZjdOYfI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qfQO4VdbKTpU6s25roZ9u0W2IQ08y+6LFnuMKThrKN1hhqSYoKZqaxCw7+7+dOwYONUoVDh6Wi59
Y+hGQ6HVycgFcoV3PaEcdVB0RoESzqmpiYJ6SrD7h8mfEIcp8t/XKFfDABpO6nrhgegzhtWEYOGW
zNnM/aMonrPoXnt40S3FQWlio5xbBJxLFXmdWCC1wAOsQdYsVK8EQJIFPrau95y+alu7rU9ksc+/
3L14+fqyd229GgD6dpTKDZDDB4x9rEW8XXVQwPX0lSPpwjPUyfMNaFv3y5Qs5okbJBAUJO+a4OxB
UKx1FvIAwLTAhlwqHDdnjdWxezTwyvyk0LCzug==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tm5E70kopcZVk2lyLZL2DhsNkZZ9007bUVlLF0bQzFHvYXYgcsXAQwflg5D1YrTQxGemPecou1PI
Wg3CmGsY5A9b6uGz1Xjtt6J/eMcflQGIF0plxkFJ9Yh0+Ud7+r8n4mljCP6SGYZHkRKF7XmNsEdo
vHkHZqPf2LZqnoTfmz875NP1mZsee1CGNEDbbZ1ILj8vkJo1u8ENiebnBG6kJtocnIpotFSnXK61
5FL1/B4oI0S4Us4bs5vvGLigC1RPIv1QZ9y0LcCax4QWJvscGfW/bGdGhqFZXQpbYuMzfxl6GI6w
wh7v2MHjv+Lr2OrwkHgkZx+XLyAwfzJL/FyEKA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wpqBV3cdN1DAgn0KCpa1kC9lWQ1VJzcuAx5h8HQTGLCAzRUFQnCa/EFt6R0Qy7R3hEJGwHtvMUHP
h5h22kDwO5bAhKqaf1yU2gCwDqXG3DewDm2wwPj3TBQ5BBHJapwykdeKGMkQImwpxaRWQvu6I3xK
IUFYyggVvKKZnjDCYJHQIqubpmbB3Z3L3Z7uiKTwmQU0S5eCklRLzKPcMiaVKsrXf/3wA9mLjywg
udEIgv3oufyZDG+pbbDReiiG46DHu4cKmfKmIhwVc68tb/KLSnrROnfM1e43PKLLlC2Nb57FzIFr
D0AvLBs1wTe5j0nEI6Po55dq7Mi3efdkT/iW2w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 96624)
`protect data_block
CMjNT9ycdQMrEYHxTUBCKU9Pjh9de9rR2Usa0ik1GvrQ7GY0KeRrr75ksREU5zkmulB4I7/CGUIx
/O6MBZueN9/X5F+25olUPZTSfEYGtny/uV379QXZqVncY4HJRwxTcLNMqSs+aoXxptQJfqey0zwR
Qx/qjldAuM9lHvix1Ol8UPcnLqePwJm5Xp64o7Y2DJpy8B06z4YTic7Paj1s3qXNoC76rmHFXAj/
gL0Y5MV8HiW6jeX2EN1+qYgmAFWaF9qJcA7B6Ot8+pNRd4t2CkeaAqwb/Vx95Q7+Tc8mmhg/AKn9
rOz9IT8Zj+EY2WIglvSphQt9lItq1R/HA433bBRNL3qlG7/fmPRMoLpnROyraArW1rLXnJQsMDXP
Q2m+ofznQtVVQnvzjMbCzonaH2PfiLTXtVe9p51YHi11ih7d7GUYB4tlijWFTPUKF+DhmHD/thWO
+lk/4CXBRtblYn72ZABoRhbce9Q7o+uLzdz8aJYhbRRFfLm6cweHkatU8ocTG+Hbd8M9oUT7PkUQ
fjNrpvoOOAs6G1Uymzq6nIV8Yd8I2HEDz4VYFCPPVX1W8T0GHIBVcEp+C+6myoAtPiVOggiPPK1u
kdEZkRTbytIxF3QA6fvsV6Qjw6gMqudt06hetk9HMQEq7w0poi5q/lGrlyrvcYTuv1zHyGK1zEgR
yOPMCEtbzgOws/rGig/NvP+aS2S4EuwV74N/oqzWVPFZvoia6ZrUfn1eKX1tOlyi7ehFBkv4Tb8l
8C/WCwwjZijXPnUqPISzoiLJp/7SbYBQpm1+rY2lnWT0EGYjEc/itjoZKOOfXOogZ5NcOdH5YxFH
l56tdndV+m5mvh3LIzewgd+s32644aV1UCofoV53dSvZyheEydPWPHdWIPoa9xfBADTR7aUT5+zY
LsL4RPnyBpCJPW3lV1b/bUgKzOI7XXQJ5D7n27OvHHv8zvcGsVx/5WX4vhBGuNeCoDnhqr2O+HCV
7/78BdZtTgOKMYjkj2eMzilfVLpskWrYN2CUf/YwAk4foGMYUTcvY6wl+VyjIMNYxiNG7JyDkSuU
UKkBXvKsvhwbksR6ypZHGXVf8BG9vCO3ehOy1sdqgprpeZfGrlrV6gsDY9oqVSSX0WLQ4hjuNipm
E3ADbFmB2QgfJe1QSmRJpiYwDTVjKImPPwnQfDEgaoIDQQaP3HLSocPCN/oG9CoNlfEmELgmzsma
NN1XzqXdsvdXJjTtIoSDyqdCbZEGZ5qv4+FS2TZ+cb5EAhnok93470siIYRAWPHZ7KvIrykkTjyc
lRe71KtpQmnFNaLiDW6zlho16rCNE4wrTaJyL6PgK0SveiLYxFJDnDYGMqMbcO3WAhKAfTO/CQPS
Egf+TAR4UDCQv5B1euGiu9vaWxZunRnBSkKN0VTUH5PEQ99/J0h3nToeBbJV93/tHrxyL0qZMUSs
eHRPbD+B46mzFAhqlTrpgbukhhZsY5ptawTKlQFOwasq9TqFmz64bUoTxKWkC+/zh86wtottGURU
loDUPpomhlSo+LV0RzPjnpaudQKOrCMrwjPAobzK6HuNpjGrL/nhWQgmCBeWR4IWvoOtPZLMpOft
UTjcUcPOlVJT97jzWLqgPlt1o4plUVP9noZ26n/CpWHmkfor3Mu/qs+SVnROF+ZRvhAbrwe8afyY
JacBs1CK+vgE8Fouqk9llGWG+/fanotGG7jDLkZ8ZEC3dQym+Kkp8ybLodk9yUDC1R0SW0fD5DDv
Gys1OLIHw8jfNpB6+ZhvaDmUEJDeC7ecGMWS5Jklnp2fWIe+tUftB/AN73vkSaMl5Ee5Yn4sFUbr
pgBoVMLiTz+a2hDEzKYNO/KDDpbyS4HGNnsAPM6cZoEvQGfZYncuF4SQWpVPsWzo2NJ+0oroC+0n
85fEwzlmMKySg4IiAlpgVGQxkfJtwPx7OhEJ61uvyKXUM148FX/Qd0MBvME0oQcidWasJegyhBw7
7iZQvcQqKdz2+XjiFcftTFwG6WzAoyDplDKHnr6UEOXy85Up89wpZPG9G6/5BdpRD4PnS5PPZIHf
kn9vw5aAK/WWNBfuH5637GyWafg61UIvlENVdRvY64zrqHWzAoxMjmEhZeMl206EyJCkpVvsxkdM
98bhP2c3j+TyEJh3FbSZNFPLDyz6gc3W0OmQ1LBzaY4LxhVMc4tVd5tDr7/pydHgFhYR96gCSU/n
zIgga08h8e62p7DAkJqWXkXTQKDpR3/Gikh9Z9sLROXkjTj26IYbHuykCo1w2RrioMe5O27DucPj
YMUxOJAMvKqUw46SLJeH6XqEixrfTrzxNw0pYBJ2NV1Q+prGNaQQwzSlc789O/HyseR9hjOOgRJF
2HmRLwKf6w4ntYv3/ir0mhyg69mm27A0BpCC/IXt7IRmPzuzc/e6X3bMiGShKY7LMFtrpTwoxi18
BEZNTfmlfqUkkj4VIAYKZs4HBW0Bfra4F9EN/TNnybgDgVm5ODihsygLV2AlgTFbHqxA15Z0EF0t
lGxxu6dHJd89f+HkUerD/l2nspzPZvnblexedY/UY1GXJq5+NtDpPYi1Eq9/Iv9YS01Bwhybu4z7
pEFr+slSEsgDwZJze6xpyvzZMCxTcAJyMAL55IA4FYh4lJ84v753HCcktJ9/NwPMOAaU34iinnSj
XhUkFQanXyxPoGvj8OBSSulxRWwGvqsLvZWvt6KFa8RtiZbBeEQRuLo7f1axGHR3LsZj/FPEL6s5
1aPn81bt1SIILwP4BLD0xoSE3sC6Jg/enr/WqMjz7l2l6lPJRh+H3K2Ow06ZZtNRiz2xaVYqBPtr
C0LrqODRPbzIv96d+KnG9AZ7y7yPBszXIZiHaarjR8ok3CAgQnRQhJ5RfmMwBthPAU1X3/cHV0EP
NQHk2oS3E6aF6ybFuAaz4XYqAaB5CXIN57vjwaUg1NdisVapt4eenn7FWy3495QTKA+8YGNp4sOv
nyrx+E+wMGNO0el/84iRbkfeDY2u+nj6HHCt8CYz4552AFzcNcJIGwVwfjsEvTVoDHzTw3cBKBam
9GyLMvTdEj8edj1oBwhM3B4i10weaWGdk1bcmZvAbQtJ4hgzfCFtVBe1+rrTm1UgEfSJqlHJ+GMk
gi7Vba2QgzA9cDP6OWW8g3P/zMf/gwRpuNuJdLiYNH0pDvJwkSzuV0HiMX7lvckCKA2OsKsxZuuN
1eaAPoLpFKPr7vNTqs92lHACqwIP6jNOtkG9yi5tLvuuRms7wXsjAUXpI/35jeAJcET7PJr0OGy0
+cch1jxekLw1PytmjFGbjtc6oAegSwZc0AIkNxXZlWcjseE5Vx0yEwuCTo5dwVs9IkCHYUD+j7UW
81EeGqhymeYtnwnl5VZRsrtkyhR1taMYRARTi+2RGai86fu4DhPmchvR/+695WWnA/JPgFQwmJwq
0wajo9vToNSPTkea0h3/Wi4+8R9CpwKc1HOTDptCZxdtT0i5D+BuEO9ZiEYrUwLyYlksUDK9BQx9
LBUQNMYsIYi69M6K8bF1uXZhnu88wjZ7i7WpsWTu3rTDhWSMii7JsuT9QoF9KUa0Zp+MD1S2DkSk
qto3k+NDy+vxIfVy70mgHB/RStOVU4OtZsyOo0gU73lV2g2ORW6Aw/jI69NSQgPNkOrvePnafn1V
ipKPS0RMWXE6RMhgWDS8dkZdLjfhEjiCbE+1gcPL3OJsVe8/B8Omm29aEFzsVCVEoPmrUXGBOVK2
eqiYCA4jctvHdT5oN+YnQWUujTYCqOeWDOPviNw1jCE/u4bUVwoLNKHngZ8GTzAHvDd1FqeSbc2F
cSTKNX3bX/Hp6slt8LphI3YfQ+0EXtNHVZ/FWAxgQsolm0jfEZCo9CjGFwWOywplHngK30smiGoB
V8iBxaJ9E36qyeJNTf59HifoNSu0RYAd/2Ru09tz+GXlaCtBIpb7Lhq2S4FoSBVJIP/JZgxkvP9Z
udXz/y8q2BUV0VH38xdjmwWx0PLiTN2ICDUZobSMzFyKyzmAHP7FnhS9fLqDMtClFrOo0EgOp4US
cxpDg5aN4imSk9P40bPC86hnWZdFtOW3qtEYuLXHPSYkLJK6KnbmZWsj+IRIdhDy1Iq8sA2fsZ2t
aEk7cZaRJTys/vw9zpoAt5vUiqX/eG5x0hjidxzqQumQKxEsPDaQsNGl4VMykQq95tNstKp9CP3/
WFf1Sy83Cau/VKVwps/cK4c79FcAwkoMuEhz8ufqyRA9nldCvGK3teupcK99a4s7BmCKh6HcPL+x
0oq9HHEmqL9OP0shD3NK4tO2QMFceBpAJPeCSKzlccyZy8V7Hc5VC8RL4Au0BBVbdZO4rff/MUKs
4NOmKldXkNlfgbW/7leGlyJMuIZvS+v6qj6cCvU/+ZmdxNHcHa+u9Q7LHf3FHgLMfJVhUk5Xq9kv
QKL+wNajJLQQaF24JKNPAvgRWMakf4hreKr0k5+NPrVk5mbP/IoAWc7t3YTWhKIuInt5wRZ9O5yY
6Ofm0RCPOnj9+25MQPm1Lp9RSl0mZBy8hXX5Xa6bRsTU7OpyMgYCDGXJalPH4DP80/4cBnUjgn6W
s4KwwVnt1BcvYidEF0Tyezb5S6ia4dSXA0+JLaa/Re6x7HnTjwoMFbaYtuRGAQkI2UhNuoJwMQJ+
O2a74kvPzyUuuvi8sJlFnvVeCmCdKi+mdyoH3xi/Z6+/xHNH1aq3YFN+vU3Lrzwp6yCvEVOWLlvT
KwCjmFm6V8MU0J0kJCcHtI66cCY5RGLZEyTl7YJe+GoQpYC93ziPrmkOXNqfhf2vqpMvbKdmbzdv
bqE+ZF4FPrtpPr0CeaYjWStezGjirv/2MNanh8yvNw9zfOzjwXcWqe4B2oK4QTwvZTtGhiEevkzr
nCOA7sX9fwYe9N51xn6A4lVSBRtyFIr46uf1CVyBuPxnYHK83rfCH3n2my+B/ohEAT31HZqUGmty
L8BxeC5Sozxt0IZi4+yiCzmjv5J8SjRooE/5GwLYgDOGcRFSy0IDI8zxbqFmErZW8/BNvDqLFqDG
K+ck0QLUuZMAkELIv2hGvpdmlwDkDxzEp2UVL2g/YKxoavwrMyblpP0fb07nalBhK17VNhWWss/Z
QLLohq35zauMxt6BPnWlhW8xkoL+OOyZ9b5XLmjf7eJeDlZaa3YeSluIYU1NdxlXYANb17ksymaY
607Vznv1v1YbfmN0+cBMjkKRc40cJtfonz57qdDBuTsFkPaCxcDIym76HBntYr4W5sD93oLp6wG6
YhzMnSvUbPUX9uvieYLaw1KC4LId57qKgf9QD+1UxwswYj98QKqsAeHOuv9qYLDwpHNLx1JF4PWD
TxvmsZ5jco/RvCnMAjAvizaBFuFy6k6MVHdMf9WxHyZBHDRA92U6BmRzMP1s6crpydgjTd3SV0PL
FEeVdUbtCR+/P8Eb5rHxd9+Uv4raaV6VkC7tTPN432S0n2DY827sRo8DA8sY/sRbr9qweeXGMcS2
yxdSbj5kzlbuk2yZnMiXOL1Lsv1014eLRhfILY1oJ5MEsJlIwsNv2wcJOZx+ITGM91Awx0yt6TNr
Yojkg1vGaNOmxDw/BJZiwwNatpnn5c/uy8GiatR90L4EYic2zQA0Qeh1FY6esdQiaMkcwABOafk1
kg9ge4J4MB6U8pgM0pFLwdTb5HTuRq32E2a2ALm0NaQsLmeDM8nDnehGfiNJfYcGlHIcr81b8h8R
Pn0JVUfR9wQjYcMgg/8slfZJl9ynZK9TpokhdV0MgvXkYsnm6TteJ2Y2LDKkLKKiOZrQ57SofhIg
PnuA9Xb90ydcXSTCCit/7btKTDl33ixM7olSNac/JMVXY/WapySbOxkDqRMIzKe7S9Ums+MUSbDd
oRvELvNtl+hK9Gm0dIsCij19AZ7eiJl2yRZ0VP9athga7z11P5XsUt+q3Ml8Wu6bMmL0LFody+pc
HGC9uut1sQ+fSfFiUCC2CY5hihRk1H+KnxFlNpUlSeO/rQNLOEQeCauOaLV+yZbnMhpNy9WXBIEH
HBBHl5OBmmEGdl0TtqAdTyXGSZzyQeGx48+dilo8zFrFhMFP04Q9+1jVqtR8rbJrIave3dOFQEPe
Zg1RaOSNrRk8lJDJUw5sKTcJGBrH5s7t7ZsEu72L+EqxzlG0p3GkbUYSDrvjvUZf/zIWDau7zMlx
QTFv3fgeapuWKn1acuqEAwYoPB1SUqsfXH46UZVndE4i0N46jAW7CGWV0y2+ecG8EdqqqUVbSX2l
JynpAeLhkK1kKVl6zchPVSUustI/TDkqtdF7zPgwORtUvv41INvCQU9KvnIUmfZyaJcJo96U89pP
6r7ZAuWdFPYfkkhSB3iexJuAIb8PIyV5SS1b+2HJu71d6QTY/4oIFXGlsLC79u647+nm3EKUAoC2
BA868tKeWuW7avPcvQUdGySFYCb2GrWl8Pya71nWMza3oc9pfxf93CIK+Pnb3AuQevo3ehh02BsH
hncBnB7BtbAZuCQVp6PCklHv6mx71K6yUwl9V8IBuoOla2q0w659LEDTi6zQxqMpqsLEgilJhQfv
avZlZ6YgSovU7awT6aycAeRpzQgXIkd0P8Ia7HZwl4mYsT40mZHAdDPApgujjbVAyBSN6hQiN5i5
dT0Xajx02SifbKs5mMDwoUhilCPNL2LcQUDWsYP68Hk0JRuFOQooIrsuwEeoqU3PPLFfJ3RgU/tA
P4qPtaltNxjZYtcIBI0ZbiqNjOvUVds4xekmrGN95Pekk4feE2NgPU+mrNiDalN7P0fCtg0uUrsD
Li/3bbcTU15QtawHLEeMNJpK/+JLrzqEpeEGjLJqXvpb3/sbifRTgP8RV1YldtO0mjjvX+T+rs0c
7GWke6gFCtc2Ncy/FHqcGBzbPzJPIBarx802M+Ha2kCelf5VoR1ozhe8SrFvIGmlEdCjiF/OV6v8
C6Ub5t3rEcWpJ8TYWMydk4dyMYhH+Or2J+Vyn+asBamGWh1vsxhXCs2/3M4ip/TGyYhT90zVCSjT
WlA4sYgEiEMHOpWNnzLb9ZQEMt8066fYFLCAlxVMHEi+dBuM8BO55s/USdZFl98pL8h9HI3A8/t5
AD90p83Nf9khEB+TTK1p41Ar6TFv1zcwxmmQjic5BStNbpFP1LROzgaRda72rUixG0VBsQ1A8ACr
xxai2mC2IQ9Q6pZtMw9fQstrHI1ZrZDkTvttvELDWrTY3nSCX9rs5A5agbGug0Y4SpZcxOKyQutf
my7l1a/kjzHteLsqzvnDEt/rNotftfxv6jwrfe7aX36xMohbmHh2GveinjAYptPyjItSJXvdwLq+
gg4DxaCAKEgFQiuMMa8/caijuhojwuBSM3hGHqJZi6FoILSo/QVo8kLYUmXGZ0aFoSMgV5cN6vkC
ZJO7ByJF9j8UepiCqW4gotlZbkU8A0woZOsUTuitBm43ZauEXdPDSf8uYJ2WZvm+LNtOrNQvpUtJ
d1Hl5f72rumqTq0CES9LMDjkbJUmU27QloJyWcPtoS1kovj850rh/SJOoxvVl0PEqKGtD7cUYjSA
cErceOIDheuZP7d8CndwvXCDMD/McltxDUWGUT6km2sVh3iLXnNF5WyUcej5kFuBDbizTxgltdlq
Nun7TgHTMrkpBl/5TaTJn4fuCFn33V8KPczFVu8kj86u7NfSS5f3L2sa9yM+2jYdXGIbgN4CNKBy
ouBSDMnnQ6phif/QOvSrJPcbvEmpZi54gHjIR2cZEpR7dI78KHs7AySYq5W89BiGk/h56SUcU/U+
Oh0njME0PdtdHBwqWgP19pACxRzr1U86ZCYMCA5alLTt3hCZTMrEgj5FmkamtH5kp6usLYK8dOz9
7jf1xnyjwQ+mottvQCcWUOameU088CUiT8Uur9Dr9rjw69DUlEONstenG1wVq36l871iLGSzokvI
hF6VJ7NPtqV64/PLSD+xXsMx4JjDJN8lSINxFuHXOuAxheSGvjv+4Lu1xbTcYj1noQu85AB1MjH6
hOx5EVI8lCt3PG2RqzNpBofcEXK8buVBsfJrMKM2f7n4l7vqFjbI56S87yqw46Fu18hVgm6/yheE
5wDzAFrp4zK7GCHOBGmhqWm4hcsjvTP7BSSFtGR/6mE2nIx60dJaCWJJ8OItH8liUkt4NcUIn3zb
wWgfDU7rKUJ7/KuhkqzBsihzHmoN8bCTwWMa5IR+++CYsrpXeysHKWWUdCYsJaVTVHHLw70m1+mu
gRVDmYLxn5y6WdjmymVL2hdRTd3AJZfwCyCwbwKdjpP5xLTLUm2WBHjyn0Ld0fWJhc4LORi/34DJ
AxTsAPBXxFCl9ZBEah308yen9aqfjOIlc266CwhRyJHzgWxKxzwRrLTdiJRiXPUtjF00M8k3nw6I
GFE4CY3A7Lh2oQVWtHd0XG2mANGAPAvcPJKTiDCG3IunuD6I96EEpCwpK6hL6GqgeBVwi0P1LH6l
v15KoScJ5y2knV/Jb+Munkw2RUNUOWP8vXgNxPphRis0d+kJn5KGkdBA20ui9TeVsp1B6cijwU6J
Fi7iZhhw8wKlgzEQWl13dpV7SFZCrsJrx4khl6FTQyQ93x0ONYUMhOxk+TFX4TnXpYH1C8SDdHyE
1shoSthmv8xVeRrhm65uzX57+7x+zTl4XtDBIomRQyWndx7IskmJAEZCmzlogR3/5cwmns45D5Du
MD9drkqWAoVfZttGqJTfCFgHgkLOB5FC2+/qEUSNKOyEP42JBomcBdWxJexKE1Cbb9SQC+COWhCp
g4UorlVNzK6JxB1d6TcviVUNWonevTYf9/6S7BheJRU/1WJ/9YC8yd8BP0eAHO4eCO20/lpXLlwP
sQQ9uhMrREWncXyoCClcLk56X2YZRGFU3g21tflIMmc8H03/VplWLctsXWyTeHJOHuLi9fLfxnzr
mgUFy8ofbe0yDYAeCulRKwVYttCpccFwkUw8J2AxeGOidX6iZnu+k7XgkzEp6/DNK6taYQdNOVSd
NpN74GUGmzw4au3KUSGMSF5Nhze+815pBpT0jE6ZwvUscPFwrC0vFLyE1W54cVYopxje+BgBOR31
6Ly7sVwzgqtuNO3UX+axAkhH5bokWkqurdqTtyqqu/W7+acBSAYxiGKLd0rYZc0+khKEnW/FCKbx
x2bwldhxI4jRsOSfwSbPVIeDKy67zdEnUXOTgg92iIAEzSK3UNBlSSwGaHgpnLRLiJypTnd3oPmV
HbWtoZkwCu7rzHOC5CG7WG5IVLNjsbOfFfKbdCoaQ1tj/L0l1W/ZmsPA0L7vYCY0KcXG0lFzifTj
jjD6A2erTBHpqAe5vGWL11YEmO6yQQHmL+6NBLGy6eC+oY3nvaAKDh3xwon0mSNEPQX7aQfAdFn9
bmPsscnApswCoMH2zO7oAlGftT1AotWtp36KR1Hof/tZpY/+fA4a0hDm0oFZgFEuFFExxCuY45st
4j113mG7PPAWrhvaFji+EqlaAQ6SRsAQ8UC4mrfqcLnW1Xb/bypj3XPMgmS+FOG8p6xm7gJRW2rT
VGKg4SspB/r82gT3L1abUKwTTT0QWuKBl+tesDU4LxZd7Ee2nVLqPQ38d4JlyIGxMo7vUVQjTSlY
sayOh7Tynjupbrq8azpG0hvMsYB86ZyyOgAOHZZ4iBJeW1ThaR/sru4il2u4owA3sKq3JbpuFsDi
+JEhbd7QtjwjebZ2hPrqyHK7dUn5GEsLDZWJduT6eMI+7AUHwHMCAsZbNA57OyXdRcqaw/cw2KT3
/ScQ7rIc+flJBiWdgVRjc9WqEEudTufDmXdClCeDUdYTIxLtPl6LiEzjMlt0HObbJtLiiL8NJnSc
oP9imCvjY06gGtXQdBmAn9t+MnRUUW3XqLnwe4n3ZANH669HVLqmokx7n2A0N8RfylhQ7Av7apOp
ycipdHUPFdikODXaw2DSPc97yAFXGMmOZmUJ0Tv8NgXBDsG22fL4iw2vr2KUQ4pfl8DrVMC5frJO
ofsTZPM7C/rqLbeCiP2y0TCOGVDe7by4slQMr6PXY+zOPwmBlETDIASAI75RYCNPR8ZJvcMRpr+i
79tWMKrOmWHoZ032RXxUiUHmpARrf9zuKfURlHLWlsvzyD31K2WVtsmB+NxkmS/c4vQgCviaMoK1
rwpbuudZwSls1ztldIt46Cay6Ry0lRWky2dcvxwTnKH3uiJcblM3u9htK2L0VHNo4q/3oe8a9Qys
kz2chnqNLsct3OFig3Ps65O2SUS+p+2GdJ7eKkbcXgm8QF29m2sMzHymoz4ZMk380wkzrjnAbwcz
tvfLu8AR3LzAebzwh69z4zuxeM3I84tL+Lmt4HEibdot93/AghqkbZDOUsVZer4+aken9OFeLSUo
seCR0GHREP/eSOvXdh2OVlEozNSn5PKzgzJQk+mJqGL0+qkeShmXInq0bMk9dyR6Fy9oku27yc0y
z2F/gMhn+ErKB/VOcTcSmIkRtJXL4xG52LfwBnrQOnwo6cdkMqL301ZobUTpw2lLpFehOPCeplm4
/wdDkDjVVrzRRFU1tjuxoVDrsV1yNPQbH0V5cXw9sXCrw76F+1xshn1JWXKiFStSyCHTuC2WxkEy
WmMhaVyKS03ukfXW4v5+VGzBw/4KiPbH08+LFRhjAzC0bnjAhUyUvERWkZQeQF1qQYWGJA+ARY0c
OeuL6cWWekzJk0uRWMniU4uY5OrUOB/J7DlC2kTvVWu790pYBfe1dJOaKUOxIS1e7ep+6HAdxfVH
Ayy6DAgAIBtUxzB8hES9EDZ5GPUWUR1+T4Y+xg/O4nW6fDEi3wcyPEvz767CuaDxKJ2QjhTQjO/P
F2i8TWA1WXJRjarQvgXHkiqyGEHZxsO9xX5Dw6xm3NlUo3vKEkrcjyuJjlm6F/0Xv/je5LnC+SHp
XYUOMNiYwPgPN1ABgBaodiKf/9L7YSGs3kSRCTJF6c78HbRk2css3OaEpwzQPcb9IagnSpK25SFC
uWQjHuokxiHLA73bk1RKAnauRE/r7ty+0Ccq66LrudZFV6DEpGTmAS4B8bhMM62JmP9+RuuxAp9H
qh16yZmeNuGnhIkKMkSZnIlmNvCQ9Dxf4CRqOKnaFkZdsAIRxRL6KISzX3mC446TGJhtgwHHBJeP
TBTBbHcAaQS+fXyPFdsya1UoW+9+2c0y4bAE3r4CqYLgkA7lm1ZB6HTRC1p2LVP+nX5H71R7+5q0
PnP/mXYxgvd36c3ZLFoY/TSR6Tmj6VCwushKic89SYX3mlMtWUGk3rtlCugyU65qlNHNI8C10FX1
zinV3dg5X7+A7C6NfB9tz1+n+FIz78xUP5wGMP8yTyrSU/8xEGpaTyO8UB4dd044LNUDfE6/wy40
9TSdaXk39zH+fSEuvu9h1FgK0S6SP+pZXsS4U6ITOBIbbME3fsxx7bnmYKGSpMuW3H6FuX2/lZz4
nFRyc+Pk92pZ4VsrXOkQwi62hVNiYkgeZdCluGKZsZ4obrZHMYA/BoVFMzebwHbj5yLzsOtFe2HS
jQYDbuuqPi+6kYuc4zFawcazocvEydb1yQKB2NfLyUwlomrSkV8HtHYieYpjq8goq+K66vJkSkCS
4Mkjt6R3fuaKqzkIpVdN7zPyHuE/155aNB7hkMrH/V46At/YZ8FzhOGzBx0r2ru528/gCFqBmKZd
h8hw70MdK75f52FsXs2rg/4B9/43HXvQ1i6laNJjOjAjyBo92Ndco2/YR8DsIZ9Poalc4NIRPxVG
ix8PCqHpb/5NyYMrtflLv3dS9my0k+7fUwXkuN+TGpudpxrUrloHhpiiCr+jwzA6gdQ05EZnbcuO
jZcGJ7VJDUjnAm+87PuNla7O2yuKoxLP7LsD5NtIC9k4cHpZDu3k9/7k6GKoZBOvxOYTIgNhhNVF
RfWKzuFnqcUoxXRpfG5NflOf+surJKeimwwoE/UZMMdfiyDWGsdhN1CCUMKIOPKZ7DIjz1+GAuxd
H0/ZBRimjnqAtia0OqSgsEI+k+0qk/cCFmRSjojapRotOPDj+or6LdLnn5sq5Oh/wAQo6GVe0+da
9NUMn+9Ebg5sdrcXdjbOrWRjBCK4A9vBfHz6o7L/cWGdimIt1P04dimJSQt/JiImoJ//bYVSXFQx
yWtbWkYLtwJwAUY1Uqihh7ZoIGIybrgH9ysUrrOaHLtRcbLJHw4Bl6tA7PdLMm1H/LGCk7QdFHgQ
Iqz4OdIYdTfp6i3yZTZymHzxq9aYblv1KG1VjGuVuDRPvH2kMS9AjirGofQUWEpWKeKwW31SckcI
FVFNhL87GXqup54HX+IS2fJyxfzCR7f+EcyUiTbIDNv5oWFoYa0Eca8E8W/eUQZxZut3+4Ik6+4A
eaAK1Qm7josgSjcEcN4hzOJ7AyrVGvdWUj2qg3+W381xwtSJVilVByN8wroCxABeB6PKa0Mwb3Vv
+eLKRXluC9pgM4dcghdKkx5JwtypHdQWr4PsyDc/3lcFVPiaORJyZBPM2adoU74Jv0IS8XHjvQtl
qAt0NMjwVbQpRj7WfR2zipjXuB9nwuVF9krUXd+jvcL7QpdjK6R2bcAGBx4uMJxJcYPRW5UU6Gfw
YZ2sSqUycChmn81fSKM3e3CkxHJtGi7CdAvL+Ivok9d5jka4chAqphladhvhbyu5qDdKDujfAOnB
jV1EtzNOWiu2BOY7dBpZqHN6QJoBAPTeSgx/IHv7Q3OM14zPiQTKFyyLw6BfnMq1e9X23pTXBHJJ
4Vm3BbqqvLtdmO8oW9X6XwQ7m4pKnVhfKdtit6oj8EGQHLmkE+N63NFvHd7xiu0psnN1ZBxeV538
xiihkeCtZl/BWsu0TfZLX4ReITRBPh+OPFV/IW7tl0CNVkp3uTfiW9L0W+Q8sP6Op6clcYsMXjuz
npp9kCuCcOvUZaPhmTucNNFQcLNxpGIY6A5z3aGJY1/UOd7cG5hiFbbE62oDOo9OipR8HDgm4OYf
ObedEHLnJCX9+Ln/EmXBoZ2N4raCz1Hk9Uoa7L70SiBAce2AzC0EcCeZHmsiac06O8lZv7ly8aqJ
z2MsQYeVTokx8at5ZFxw16rJR1jY9kxm+ZulxFA2Uiv5pFOuy4gtesUfr2J/AYNao3qsu9OjARCe
f52LwTXaGF/VXBBAYkRfi/vOd7650PIwYtmCa1/65FhromCnaCUyEun46/wAsreFAXfrjL5cpT8r
aOXeBO1Rg7fNWUDJmUP2s4Csu4+KlpVS0gH+fYv0AzReKLNgkBCtsAr+WyjUGLrzjsLCZyCuugrl
4kPXGCIj/8SoBGrcJosAyaO3WhRm8L0PrXWyEvn2oNr5XO4FjHrgzsQHDhY9V51o8GldOH1MD1Mu
9uLUlCXfAkQUzFl/Twt6KDCwvr3RTtfDOuUbkPP72bbzFUv6o9AGoD3ayq4c26JP2kRnGpQKfWPE
/nKa8njQdv3Av9lOxCHDsRNxxXJ+UImDdVa3TyAPnDQyFDmg0ybr4iTTQmYUSbx+5brwiyf7DjuP
vmD3zCl5ZGCbVS9tz9Z0yN1rj1ZPmATu/M/8E4IihEnZT/3cbZZH3X24iWyHHTz6//qXNYPE9J+d
jE75GMTixJEqNNTt2jVr8/V7AUsPdk8pB9Hf9HrrfjeYjVaNcJ/4xZjTzwzqwZvVQYG5M77gNcdn
41Tnu7kcDzggtfnxRO/eKu6XW5kh2zXYY1QfraVdtbfv9gom0VDDGTRkLTzH8vdIS+rVLIlWsAmc
Td7GTsEu8hGTUVJu2cmfL5uCMsnDm9MrhUS5J2Gp10qNi7FdqNsISgZCf2LOVjNLrfdZYSqIzEY7
Z0lkiHr5+COBSqzaTm1xS2nhrpgNDOjGARB1VHb4CSGFzsiGhrRT95edovfHviY7O8exkwL1umNX
teBiIAXZ8FaY1XiKVEAl+wGlFh5cDj4ikO2KNWeGfI8d55laa5eaV9X9FBJx7WKTtTcEK42BeIQ9
poseArGzs2OIHllUPT48tHH+xVVdLdHSJBG1Ku8KNf4LmxaltS/5vPyv2O8hIL4pKv2MS6EF2lnk
bEYQPIJ69YUY6V3ES8uLI9nWDeWpFkqLb/wmx+F2oRATdtWgfE4y5uZYRbRPhTRaKz1t/yhw/ZWq
l3T5Nk2DFZvdwiYjnwB+MtS/cgnTA8q733B1jxRw8Ef42f9+emZ/LClpiZuYzLUrctNt6Rrw0QjL
kPbHYIbFZ+kphI6L1R7F1ySnH059hPPWzv3dBMPzvLJc/v2sklTzncZyxTwg2PXx0nQISNadyFZ8
dzZoK9MZM/6yOXvbkTccMj4uqUfRGavVQGfjaJxwvwxVrTkuoEERrR1TDjIIt1uQ32F4svDBdqzK
9ioVOncodhPya1FPznMKuRfWyNX6LZX5vgfD0Nxwd84L0z8ZD/Jnsy5UoilFzsBii8dxqqdt6JQW
OCi/Q3wma9XAu9hSGZRbWUBs6loGjV/CK8hsU0USd1r1l/PJe4aUouy/HAAn4nLDRqIqLBLXYuEJ
FpWgLqAaTuuudO7JsNwtCyw+ZJ5hjuPeXN5IEV0NqLwyrXtXbu2eRchN0DUloecvyp+lkqoa7yvk
por6JKMvLmm8oJE5AfRxDjK5AekqpjtvQaLiNqE1kPk7Kf2+lEQZ3hzI97G+bAFonVp6WSnB/jBL
zalFOH0ZtEsjkMUNy9p+NqqvScpVa8rfjG3M0MBnmNCaoqPlW3vUQpTQYZuOJt35DMIhxq9JFrlf
eLcExjmKuvKG7bfqCFcO9kySAPlSkOvljsD4uDn19eKaDH0e3Ky7dQzV6Y98GpFDPJ5aLG2+AH/1
yTora3D6yqPXsw2IWSWDj+S1vQNrPkyKyGb6iRHD5equXuP/+90Xv4SNisSBNNbHs/ffwUdr5PJ9
5CAVSr+znEK2F0RVZtDncHAlah2uNy/Ejuwsxmx9kPnE72ZJqtLH500Jf3ngxm3cuH1V1QHIdS08
2CEX444GJfztMk+I9dyCttkUOtf4PWKsynE6Rqq75hRnXoFIPbedRbucmlZDoOrBdYfSOz/JwBtT
QP9O1ETXr0jeIZ9yqgXgrJKCqLJK2jjwxqNGVmzidmMsCfgfRdlo3Je/8W2rr5p5KB+fVOPN3rqh
EzWfxSZelsEjIREGxx+bUBqO5irdowuv7l4DNPY4kKwexrjX5WcKJzLxUO6iV7OSg5VO/gGfpokU
+QYOjsT4hJGqXPNd1c0jDInY/1wYgtZvXb8UJi9QYRY5b9h75LoJq3NVDLb/RfihenKXTgEJglye
GB2s91Sx1mS6VYybWZHIYuJucW4wAgJq6f0cCJRL4kmW6w/aCqmDpmuRZrmv48o47WbvXJ9J+YcL
Qlsf9MZGQMCnEeqO9cFYrWuRujGnvZtiq4l+LRNwqKU5uXdFjYXveQlN9gt5m31C5VE2JtNwYPFO
9aZluZrLRet3lUWaBd7XMHKvFDgKIDwgu9Wt7A/ofUIAcJJCKRJ6PUzuNg5bRO3VwrUu6OMcdFG2
qeLg8vdZf2LlFOp+5R9o9K6026wQsnPmGI9Arr4BmccaqAZpyhPXziFWwafHoRkq6hj0tSppux5n
lUl3Yem+YJG9bn3M1BDcGI9S1jNf4vKVVBbYeCD8KZQ8GEHYCIE89tOo5mV3QbMfYeuM0GBkqktm
BdQiUW4qJLQt8e4SeRPvBX40D2kx7UDLaciq79SNDqaKMX2yUWpMVtHe9dKYkA7rcQEVdDHZXwUq
A9J7ralUQAIrkvufoNz5BXmpgwLEBxfQ/5uBnbLdkTWTjom3NMTwAUW4UfbEJEIg62PI5Gg3VHvM
svo5SuNpp5tUDL0N1SIbztP0K47AgFfkb1cQdHaaCZeaYthJRsgIYv6xqBKciaU5o39Jnz5xTsfj
bldv9iyCGclVfqgIRJ7UxQktgn7OMuuZxPPHZcesGlGnQYVkzZLOpSBR+7vA03HKdZaBjXiKjLdv
oVs1s4fU9VgkATQwSrJDD6jb/5+Hk7a14TCe/nI6v+VTu6AaReoJnY4Jx2leL+tdawPMZ7q8w5mt
FRp3XHyKKXyqkG8BqVo8arJQKZN0wpYkITv+SHdsv5vg7JkOhyPYXff7va91qUOcGk7xqyWpC6ft
174JEV3TGy3yjTHhnJP89ov4kb2y1JWeddAE6ztiUVB0Y7B9/wnfiTWeDv5iwOXVm0LRiqSgAPuo
u4rQ7AeqPWltzQYt1I5mHFLLUv6CLK7S4mS3Q8ouc/JCt46FxY6VnnscDDzKUdOgW01iAJj1q6A8
2jHTBW2KyNPdjW/T34ZuaiNrHqx1GIA4FOiceqiul9nmOekM4jrosRzi6oSA3FTO7x+EJ2qx2STD
lWOumJ/3/SXz2UWW3f3QyzoyqUm0GQ7ZTIChpVZzzYj4dtrj1cf0LkRbzjtkW7rDKfB5aDf30G02
c9O53nAlrtutU642onHxIaMuAf184tu9O9nLKUC0mi0WNRkkjCKaSCW/vf8lCkzoFRzQlmg4XHph
l60aNTK9E7qj9vGJvmm0Mzm2Fzh1KCTHiYDXTIjVb++6DwYd6PdnTu+IrfV21siIQT4iuq/zhEcl
8OYgNTWKamG0n2t9fg6Ll3+jfLBq7+GdWH0qef/BAfZUMvB35+KZK/4zyCt36NaavnGaCSrUDBdS
rOg6aV/Pmb/0NglMOv6T4WyGnJzqXg7RSpxqbVpCm9eO827KxEuj7ytoP3Sf/vMB4P0qUVIIaUF5
lgQSYY55enUKOxXnVi/fLek+AUGtsig4mZhBRMPv+DhdEgh1dXIzPakL8GnLztFlE4Rc5quc4mjb
jmLopa5V24kMnShQaCJQLQbOI9zBJATG/bLZ1jzj0Lc5qZXnX10Pdf1r//8+F1ZDyGB4vnRpL/CM
PL5HF9cjWl5CKoRBCJvRUWF2QdUkVYeS81BIqZRapDH6l2YUW7+pe0I7smSMRlgUKtB5q1d3Cgy8
IPehnQhUocKDpPdiGbpOlpAUribvUbSwOCvxWhf7FZQoD4GfGwIMwQs2dyWpDiffRWO/eSBjXtD5
7C+FcjPWOiykl40VhGKqCHn7j1wlywakmHSX2pm3w8d4XJ5OgUxSzXa30Q/NVJQ1juDQ43eVyoYY
F7jyeXNqKmJ49QKDXrVacsbwEbqVIVTV8h810peTWAW3WoXwpsnv+ZrHHEdbRDCD4dQy/Pz8sBiE
tk/3TlslL0+r59gwsVdJhWroR9ZGxXMRWg82eYwMun0NLN6lxS0A+iza4Mfq0T1SqK7sOV9/fYGp
XVh4Hj11c9Zr1/nAoNgDC+pf0hDs7MrF0OFWCf+bwSUsY2ic8i4VG783FVAM0XpBKw12bqE8PiXq
M1ADDrFRS3kDWaxFB4vVpdFrDPmHbNzJzAdG7n4k9C7or0OHqT4f4xFZL54SzhtvhEsd/BlfmBne
em68siCtnttnDmsDGnjvpzp7Op2Q9nrrhc6kGgmgXJlm36drg7DxGgu0w99qZg+E0Rff+DZwhyP5
rmeuYfSMQcyaX9IU3fxn6x4Q1wZnQl5iYmjetXtwzfFHttNqBLP+eEnD4pV6O+Q5MF6N1NRkkorh
Mae+Y5rTjtBrhGLxVHeo3Ep4Flge/T+kpsu3Yl4/Fq36BcF1s0sW5kKN17xgyji21sNPYNCS9I5d
dBzQ7/zzMXLkCErYtg26xhW9dyhrIIefE8fmRjb3G7TXdMA7noTJrIrUyUf0Sm130BHCnXGfrHK4
jkYrfmGwUNm7xVdbb4nDRJUtRPUOA5kYjLQi+vEyZBT3BOVlFuzvYUMcZeJSZwLx9qeDLiOXHndo
IRjhzmOXOiasslkwFpbANKOoC8pf9d3RhBQJF/vWPE7qg5RDK8A1/1SwW22suDdsRIjbw5LDTicj
VL3QuRnTI4iIx/05WfzkSzUxT1ikp/e4R/B+v3seeQc1FaINLJex5uOijGKvMNsCAf7TjAVgtZO2
xgBGQ5QnrwXM+V083uBSvJ20k8k2kEiOA810PAu1dx1aKXUkM0avUowVN+d0ULyFlxZgY2Q+YVRY
UCqMfOT/WjZlakKZ6cZJcuAF6MCMrUAfkLG6VlV4arpz+EH01HlJH/0msvsxGQ0KakShWq2vPegl
G2ixbYr6mbPmQN5MZ3VuBR/GcNNvmT1sj+MxsX+RqhpL5/eWGBEiHpmLospu6U/KuI6LiJqlJi79
S4FR/uUJbAyOhqNZUdtXe5lk9TC8zzltYuYDqUHaMPjRx8Sylh7y/y7cicIQ2vglwwhp0w02RoNv
JJsVOfXYz+cZcXtHXTuBt7qYi5DWWkBJhE509Ig2KzhZq2k2n4Tj8GVba4Wkx8mlpHog9rDN0aln
VAp69qR+5DOQSY+sldXbVfDitMs/UsXUFDIgpwkZr7FwXV9yVm45kFgYrU7W+yWXU9NtNVDmLRJ5
7Ha13Wa/f4RkxsnAwfLRel9tQYJBDfBKI3CYKqwak4c0mML2RN9b20SbvXkj3G310/mchSYEE1QD
SAFYE0/iJ9J9+kEUhNkyzsKfyGD/KQmlE1MXVKqipPz22uZ8Q2NcFOlOfwmhQoQTCbZO8NEcT6MM
jF/vrDNREEC0XOvCLDhcAPVQeXve4EA9mYz5KfT7sP/un4VhybYFhvUpPygFfPMVLPauu9DACcKK
LYU4t3p5uJW/LCOIDuPL9QVm25xB+5EIRehrexlBqmsxk2fesiLSl1nzsYhlN75YHxS+/CCmFZAQ
NrVsXPQGK7vZzqAJ20rvqp4ylfFObOP6z9npAchUy+3ODXesc5ie6V5SAsZX7YQoNR22dRZpthUV
IiMFdF2/RLIJ4uqKhJ1UwP+IfrB/MR7MQKqleHaN3Gzon6kAJuvxiTDQqbUfxUdAiSSmdjL2AlAV
+Ijd1yFMK807rDPebUO63SQm8RW5TlmCo7X7k+YhVCHh0qKeCXEovB1iEwqrVvfFn1p/GOZwxI/x
8nTe8yFUVwQSWyQ7zJ389RwNXMQ8JRmEi2QejSNHHQin53rLiYgX+2dueee3XAGBpwxbhsMU86Uq
ZlWB4yob5/gDRWs5VdLvI6SoFj1KevB8aQ6RWPfGGf1CZ1dI3HvjZpoTrFuM60gmUcjL0qrLU1/l
YzfeLL9VCrmM2tZ5+2y/y7Y6CCXJa4UUq+JqTq+2rDZizkhsxoq1Cxo64Co7SDEvWZvYUAOWDZ53
ZlOm448E8Y5ZTaQ15aRQ/7aKAV6riAariJ4IA79ZQXocd/gNYfQEZx+9oFyP+I0Imd1xmZVBexct
FL9iuhEMgb4pdX0klgh1Rk2wkXldzGsclDzI9+qADsR1TeMk/kro1kIm80Kw9WdgASksmHYgE/iX
A64NCV4mx8NpcYZruId8xZS4DIWldBfYSo3SUmSSpY89x/+D8iqOaaEpnChT5iWJSW9VhzNFXqHG
Qo6IZLM5aWBktDa6kTZDGrV25SdMTK9Tz9JOuvJvPkN5slZDSPkeouc6ekJtcbk8KDgf50Hkqr0j
ORQ9r6Y44sGzu4iCk7Y+s0mG1yZmuXyGgwvFJylMqTPA3vsw10R4CewQd/sWYnjjAFibjOz6148g
vhnMi3mlVFQHM2CcKinu8F6AThRSd44t88HVScrgeof8suyHljejaiY4BCCCNmxyrYNLc9GbANhd
0jDD2o7kxtQG7fdHvzr/9b1G9hW5Cpn4UQWwDkVRnlEOm1h5EUBY1wEiV/w757uOeDw07XwfTkRU
0QsrZ3WkLOQMnRhJ3HKJsKpsJz0s/fvoECunHFUXwVT6z/Qq1bGZYOYDlhDtTVh0vonuwXZiL85E
ysKHmPzzr93Lvdbj9leQldEVi4iZNtM12QENH6WSw8hbh+R/8zSC348ZH4YRhC5355fhHqrF2WP1
RIWKIsJkutBAMNW+LKhoeXiySIQoKO4ZPYm0zjaPvtMU9MLwQf+e0k0leK9SW6BQ7h3XO0je8ZLi
SMkPpRYQ8t6MT1/dtdSv2etJxIF3huFJDL+Yt8rAIUxt69ATePS5OqVwiVauwiqUJ/Wm6dYjgxVO
h9lE5kbCEPf33ynVcRMkKz9Y8uxXGp98mFdTVv+sFDz6xomTUu6iAc5VJPyCvgGhS/4/ODQd5+h0
exdKdGYKQVszSDo2C+wkgKGjLfIKChsEXaJVCdz9QCb3MOrpiZY81rmqliwuE8nr89NkH0+6mCnu
LEzCjpspnQbAx5Nw5zWnQvYjEGKPsgWS1yxXbh0SEQ+wKfW/p54waHeaktYRlxGn56yhm0gj2SD9
Wy2dfQSM3nVP8t6DJrkiCejyc3NmVMB/bickgC6eO5R0cbiB2bIo5Jex/vMDpxSQowBWPsx/NMWz
4/graGKzqC3NdiwxoT/cbJFVpVFrg8v2BiFlfelk57jV+Wvl+0sDl7lxBbFMjwXypa7l4adpR0VC
1s+UDXLRsqwkEWMMTJ9fMGd/dd27mjiCuXpimmwT0b5fFUoxIccQgqLG+jipDXAnxzlzx9uCSjAw
VdWYpXjQkJ3BZ3Urr8MoHYdjx9VNI5QrJR0+uuwQhgcOCmV6OI2BqA/Qdgo8OpFGkCKr32N1tHeA
HBfebjSYSb+9Fg6KN8OURB84eavo6tYHf1jMdQS2noIjNueC3dYv9qGzRBOX9ICzOcYj65yQZoSd
sIv1eq8RFZh6Zple8W5BGPfV8l3McI7RQOgAPOaDTVNU1HxSy78at+2AaqspLf6Yrc2dEMyqCFyE
dKn6wSzOmJ2XalDd4QePGCNMZv8oHwdU5BKrvNL59WktGrjHPBpNsxhgpKEhlS84PqeWVVUhAyUq
4cgpHAkG9VmZcZvH5wR0A7baqGxJGk+B+AyFsisPjRF1z+PVjK75AuMtUaojRYpf7PyrRXY8G5R5
ML/SZgiL1XDspe42EMkQTWvJct0HifT1c8xUvWOyVjy18QUBwq7LcI9tekxvqwwNsgzsMGyRoNPA
XdIv2Igcmg521iWxoGZWA8EFK/wjj8FRTZ28lRtFBesuZzmjd74dClMFdmid5avHFPERdPTPS14V
VYiFX5bFe8ycknUQpmD7gwlQPF1vsN9iw2jNKIs7SIdXldPLhzN1XJXZSQaca+HJ3zxXBfUaUgM+
3/w9hCq8JcnHBuP32FGAUA/xyoJwOdUEVNLPPVFzHyWClMwDHTWEUHbsPeD5JdaV/FVnz0mtpQHI
iNnBXEXwecGSA5JYeh1tOADvHgzp7/G24XKfLlhtEVYmP9Ny1dh+xJNuQjJhtgwTclf7xIpYNbk8
WgfTTLsXvXyRWXNf6rjoyd7PnVPOTHIr0r9/hRgCR1hiq38eip2vlYWQmf1OpkUgRVj6fL9IJCfB
q5albghsOPohSeimDpgBcXchoqEK/8rwDBwP5zRn/T6ssHDjd0N72eThjLjcWAugq8Q8T2x8KGDG
3thv8Z5ZxfgiNMAOxsXMng89RmovqguxelISDNrSra/84hNWzRqze0KkGS6HYEjDg2DJrrAkXnrH
+cxP/e1hLKEQwYNPEsyN4K4jo4jY23A/Bj0V+a86ljJoMaRpZ27d/PYmGc+Mw9nzJdZgsMTW9Lje
cl8dzRmXCYUVVKN6RgZsp4SdHl7GT5voBmihRszqrFHuZTpD2SK2BBazIwB+NcT1h/zyDR42x1YZ
asFKjVlmMthsxLYceIXurVPoKyuhUPW3JWYMiVe6dcHs2elf4Qm3amxKRK+XZMFGsAZoM+RsHhmv
L/snIy04xGaxUlFbsKrbQXN0UizAQ+6JcMyKuu+NFdojBQnEZipU7SS6O+UAYUl3VzUZ80g3hKDz
WJ5EfxBJMQcsuLa70SfH5Kf1MkD77p+Cz7nD9UQ+8DFH5KzSgwhC6rTbLR9YRiYPYRKL1k9yhK1e
PZ7gxGPXIzNxuDOyqRmU7xP8KUJ85P4/ib1oIqEP3hQoKUxD1VuRjAXC8qMHfJsXvQ61E3s557KL
Mx2slO3Lvt2hTgoa/BtWM5YT5jvaN8shenehPNSYLfoI3zuox4QZhX/rNRjb3XcpM4M7bDuPvX/j
YrMB+3v9Esfz0rVerOU2DiHg+XfbAFGpEJfyhTXVEFdgchcOkVyg0OAKH+0JcwxDPgvhRDA4h+aJ
oObyjszNvXH1v9JxD7SEBPnjDGyoBgJeA/gq3hKkRM8bj46I+x5itTu02MKCQ6OUmZNhZjl7W5f7
uPG0ccFqug8EqmK/Le+7mu+ovbgyn1gfZHCM3L5tlFVRzfmImwbLtf5vdeQWOdtd0T/nyFOYmI5y
B8D+lFsjvFM96I1/b+7UPaFfZv05gXdYV/CzSHAv14uBH02dELPcsMGag3/ZUnvGG3mLCoBBVGse
bq9Dn4FdLDr/wUyJCZGiGhpf7jl11/NXW3c2jhdlFVzHZ6zzyWaqyqyTpfni7ivCQrWxZVjNSRQR
m5aMl049NuOhMO0Sr02bz0x4WvAg9jN67jEbzbnnB6UEBZgculja9Wbyg4aLKvN1BbGMAynizVxp
3VV7yvW6tBcdUKe9XbaZc1gOupgbGz+p/bOnZCd0ZK9Og4l0AeqWmjtiLnDLwrz/mfEVVD4LuCl7
ZfKes9A4hfowo3oWkSh2f4ouRCePPBV9CealkZN/lJ0jXtTGAaovBMtBIH3Mx2zKQxHdZLsq1aIH
9IFZ74HloqosCEjBlqtu4G3atgQeCB7gu3REyhMAxYGwk1wN5/1wZEKrUrVAuNMFygGC4u3kQH4X
6lDAyQHl6ImDrdcwKr5yXqttntBuwbwY3wgeyY/IK5aZlx5ENZhq3ZYziuBdM0Xh65i97hQlcWPC
IihPSMhdaem7qMBC19NJ0YFWt1nq3qom4E+WtgUhrxLbJH80YoYkgwj8mfiuoSxxf5r2nEHNutd5
iH7b+DTpii7wxUl5hAY0CWoJjQ0QQ/iikKnd9Af6BVChJNrQZkav15xDu3z5vWqkNjEWcgRVfMH2
DbzuCei1rfEQHyXcsAh9FkCXQw1rYGCbN7ie1QZObIxANBLU97Y84Ic703KHx0qKleb8t2tgErhX
xzG0TazwD/En+4Lrzn5+/r2+XJV93l5F6nmQ3GxqDwoz0XHb7PN4V/b/JTxsS0+IvFa73Hf+tjCI
euGDoXf2UDQ8z1izjgklcONx/JCncdziYvOnrpvuBZXRbYtHntMuTckLwdD4go72hzIJkCDSeqXL
yK9WgefreRNa3NCvY9d2G0CGw+W72gLz8XTHdOecwc6nc1pDgJVRJk4Kpc1OAhyKsiWe+KyasdvR
8FiTk7Lg0lPJy9WsplRqTtpZn2q04X23Y5cGzOmPyiwgJgXVA+KAtKKUW3bBhtZ3tFqpn78mjhd9
0hNO0imjSpKahTZ1wsA/3Dt4cgzJYVzDWTRt/p99kx31uTe9oKHQYGNR1lZE7g5mX2RpqJiSLdGG
4I2xOMu/6yks5jvh2Dl6JPBm92cAJKvOArTk8DG3ROwNT7YwKtyCavHB+iGRxyIQqWDMp2uW8R17
c2qaw3zVGjduxZzX5LKh+kbabATwL538FdQOTmeH1k6ysXMtHvYmqnyKrvOZ6sNYI47rfVxrYtqI
kCvK6mAxCZQ8eHTIm/bIrqn0M3xsgS3pWnmOrGiN8UXSD3aQ9lKBoAmws4aCso+jhLH4RXke2asx
bqFZnADMb8NEOxJRT5E8IwZT8DuV7i5CP68XbJJyKKORNMHy8AP3iEGmue+p67zMOEHf1k0HAZNT
rj+bIAo1jTxZzxAgAR723+l+bDOiOiPCRRPpR+RQmJ6h6AetlrQbZfwDIICPSHToytyFSUE7DzXC
D9Kd3sv2tyMb/LPNtbamdBNFv3ghGJAGv/w7NUjvOxqMFmidwhGE9wLz2V5AEN8OB49rw6LuNRBy
hT6rg9FDTDcLU1J/AmX9cJR/ecVPmEavZy7T9PFC5QTA3EKdTPhAHgX3R7+mRkqjoXCscgeLgfUz
p8Wc/V1swZIsFhrfbtZC5HfUbofDy+lb5lSwHyUbCxZMEHrxGgs/xGqeRLLomYCcDRWTAdnArIS5
NOXjjw4Da0Sj5HR2PAQK8vjlQq1bAcaiXxoiaaHtSPJzPXqZefqY8IYQRY5yeSKN5YoPWgpbu534
68C/f26Q7Mcya1EgXVoehedO944c3PDg3t6UknCwQp5NIiPxnjhCEiQ0kSW34y9cWYnIRH6R3+EB
Tb4o03rfb4y2esoJsK/9pB3ii3aX3uctLuuI4n9UnSG0XU4aNOLzth9H4yiTVvsub2JzdjvMR5vY
msVW6bY/0XVjU+rdrvOTx3ZXQiORLc0eb6QULCktP9kOqG2sKqu6Kb65wDoBBeldAhCw5/IEXCwP
zeD3YoQtLE8nGKFCVN+2b0j3zuGJ3Q2Mc4PCBELEMKy3T4AFn3WniZwsEKVa0kM36m+2ul2djq2e
q+5A7+/p2EkkIQZgNP0YnPkgqBA82fQ2AOTjnn7uytz5w1fuG5v3jyNn/EuO8bbY+i9FNnIgkmMZ
5yMQ7xQl8zd0QrvpSg9OuMkwQbTAvzPxpUHeTqJmk/yzeHsVV+XprD+2Xn8xGkXSdnE3+T1AYAWj
KV1IaXz/Bx5amm01/rGM2GSjn3/I/KGxQt0LUZ/L+6JS2PuoYibcfO5wiCdc6i0eyogWV00IYLJT
9YjzguCnxQdAZTw7+9XIKqPgVBKS6QCP0CFpTjJCFEJVbnwg1vS/SlzWTz4BXGhMW+rbB5W8/l0O
VaxZDFeTarEoZ279d5dV8isR2Wt1iMPGttefUZ14yP7BYLtg9Ua6dreDHZkuVjGmh7GqnAkIizoS
D3UoXlnSSW7yPwms4LUYX4bLiAdtondQfmqg4WaWfrFYxVYUgmtrOIhvNOd6Ty9vsX1Yavv8iiIJ
7ey65FxHwr8nPwnXCrVNPWVrIUTauIuOCPO+ji1wAM0GskENeFImUeqjBXhV+65fFNJxjgpgXJLz
Z0RfQYmNlGK2fN4/z8XVpwaEUp3FYAHBzb8IFpxXGFHo1L+cCH0oL0p+UhV6uhl0OcdzkWSgdisJ
D9gC2ejs4U1/4a8nRFUCITipzUeFMbpgPgyCndhWN0Iohm0jTAjKM/3hnZDbfM1qM3kNdNkEFvAJ
lrWAIf50buqghOAdnH1eZ2rcgTXQmm7EGTLDseP0weqP64B+nRnlFAu5cArQD3R6HRvI+DSjrqpE
paHXL5o7YQ8yQjomB0AzyAkkkRXEOLZPtH3InXKVYzCoEHqEeSqa864oYM276peEOBaVmsY3nBy+
LTUSJxWc0nd48qDy8Fxmp9xwgLBOIUjNsb+BFgRWaSu2O/6kcb9bblwp6gI2HiFw+BmQB53esGjp
y4OSrptvg5HAvzXN2sf19/SyjWcDcYr10FIau1JrdAvU3O4/RZasJNOByI9j5Gx2ngKRX3rWpRHG
TtqLJl5U6wWSaCzzbQ5KrCu10eg3N+c9YRZX4vGKIp8VmSXtmjCCA2wCCNckn8byEvtrQl0uu4rI
Tr/BnJu+rFsjfGDmcZ9zHWS3suMzW1nTdZeXieeSIRNqYIo50r+w9Fz1zAF6ri4TCERApfdZZVyJ
Zz7J0zAdUvRnkUUkwoqUzactt08PUP3ADMefWvHx8l/wVamCWaATfPI+C0GIhyyby0BQo5ILpYdc
w1Ma6rNXv3H039BTWx8J3W+nwcHffsmIUC9khAo0df54eMprNA0k06d/bSaQw+BOtupAkqPs/s5u
QfGI9nnSEby3otUenUR6GEp0Z4CczYU7iVDzTzr/SLiegJ8fws+c2fuLEdE+PPFPl0uIparRl3fa
M4mgl7Q87mTGZjo0gyFuTGlIzWxfxFCjoEQ0aBBbesspEX7nRQBAzkaWgS5RwdVMwmkHqQ+/NozJ
EHt5ia6jnJt3TqaTcUPiaV40txxa5FKR7PXyAl2lLarIMSH4n36ny05SBXl0HmX9k57TkWz8HQFq
NlMIk/jbspZz1vHn0acQGj7Z/qDJsN0YB3D0U9wH/aI1to/oygOOsRCXG1YQzRSrr+6iJDeI8c16
x+O/EmV9qUYTDcTRoUtmaiP5R3MIFbpHuzaStRiVwUQIt2AejxuJRg1AQ/aXvhZLEps/uCAyri87
cwd1TrVyZi+2FugeVOgT9oIejbS0wmiztyVVUsG7UlOpLa8O7YNJpNQNvtjrgGuvcDbvO2orYI/G
GZj9JzWvlkua8Sug9ghxu1cwmdQCIOPbra/79755WO+yqMaB2vhiJ3uB258Q547ZbtEYrMeQsNKh
1XpoyDyDq5/xDAsO8uZvtKSq493nr96ENW/Gw5/xrIicyMj1+lHBVI7rr05QAnGoEt+Lcpibz7Vh
RN1AeFAOM+sQOY4BzOApsnHKMhHuqcxQfiMQzGC18qNJYAX3TX8GN0/1xXUwOcovx3cZOoFfl4lf
nyQZDEknpzXPUzj98qL6Z3C6npsSb/TKs0G6gCRiF3X79LSLmHeEJ8egnj861bIVPmfTPdVqhdPx
Ck0fUw6k3VEXXTEzwIqAj+O2mp/EwZNvjoVHo1z5JC3EA+Sr98VPjw0isJ7JhKAtZD1t+NH29Vhz
eMBX8sArXG0HZCKh7BgxInlQQ05kg4AJgqpIKjTtE447IiRZlblkeOuGlGz8wlrKM3f2l/7FUfb/
+aIuewN9XTBE7QIKkGMJVPnSlPOIEyQNYlflIQe3KZTIZ39nU9EugyhVH9txD6vk4p4VuhJtLs99
H0klVp/R9pn1nG4IK0LkKMndzNOZOy1GYKKcdkxnIOeJmD9hf+M9ZbbYxqARyHqOJOTBYevtSl0x
ZkdBSR9u1NZEnBwF7U5Cb59mqIUhvmdyySwIvYxKbmKEGjQLsZCIPzSROIUhkG4zG2mURjTd15TL
40IwPI112pcfaDyaoX9GwtR2QkA3MjgPAx/CAoyW9Ax6EEvNUyTnag35MFrazzbH4jRQ+d4HJ/jh
IElcNcQT+kx99+pQDTiLSku82Vz7+6kEn9drNWtDZaKBHfHlGqXxzwJ3N1M8TW6BTFZpy0anF46S
aUK8tpvc1vDKVvHz1DM/iGkXskWtJVZAJ1fbLtPgECkwaNu3U2l8L9wGVvIakyX3EK7gFzWXr8Gm
7MbJtRi8XuYc0+uuJtq+sIMD7+aYC8UL6pjLrJC0o4ZqHPyp6jIV+EvaqMZ3ZGBUb2fmEqwwIK+h
M2vNxHPue5CftxVxgZWR+ZvsgQrYr+5tHKvUWmovRZbGkZonrZq4i6dzR1YP+zF0ACXSQ/3EN2Or
17qzIOLSjKf6FzbD/jlC4pG+c9aWxUVZg8h87VE5IDl/tALf43HWHyqHFibteyt/BZKZEzYC/LbN
A3hvkB5xVRE8pONRzb5Sfn+lDvDnmYC8+mvaUCJQGS6/QfhwGFObaREh2/AlVwbq62vqV3tDVVml
ceURnclgWg5Y+ejiqcb6jcedYGVChdFgGId1bnayxlwo+4REFf/W5HXQrUjFVlSi2VtkgzmMbHLg
TMJ6DMUCR9yBs6bPR6xIvMMc13C0dSURAa8Q96WpdJH/oU3CggLghpdOHuNsj8SpA3pBL54eWO8z
eY9kedirQI8keD4yZ8Sb0P82qjUhXjRQ6z9qcA2ypLs9f32JmNHyi/Ez51NCl3gV48oyO4/szSzY
q7ClmduHwHapI7wnAb8O5mNEO/3I5lmrnwbTWe0zJLzLx8ZCiTsdDuyI4tmqkqXCT8zNt0zeeZrw
F5hfe41vUimVFzeUMEAFOxLAlGibJKjjLVk7h0Bcs6A4PESdKfCGyNZJCfCSvNRx5I3QKVbcyAgA
XdVymvwN/Le9VSPcjcXBtIjxp3GwYO8WqfiH4gIeB/5SP4XAuQu574J7dznh5PzoboSit6+mbKcg
OJaDg23t9TRGSjX5/Ki0iNSGOqQBKx0DcQ8rPNYnWTzzlcFM4cGTe4/kIw6W8HQFT81k5b5F1pnW
nqr7NAN2FeRuyGvATfeq1lvr6Ru1VPC6+npGjIyDY0BxuokYNr5T2rZm3aQGlAstNoiqn9FpnJb5
aF5y3q+ma3jZ93UfQS2UpfDJS50R0HtHnBxPaT+hu0StOYbZHZLQChnt2EbOqpGs9qiB0ebp/SuX
mdEwABKJrMD/QGsDX6Xd2ywOaXyc8Q2+v7SB6V90bPbfDrttL8SI2PjlLiNp4Zc/n4Qbd1sYrSgt
/rX5cgmzAJ+zYXlzJXHffkckZu3fqIgSjtsCdx0EnWk2mbWZ1dz/tlfKhyttBjd5/9aLJQus95SI
LKQBPsaS6nBOeO+hqTG+vKrdTwOwuWZQRHtvFbkNKBeRmEqgkICSqxBZBLX8TFPVXu9X/MJ8sVPj
6zJM/wsElwV7cn8xJ+bmqH811dIquU78sS8bYjNn9iDG41Ka/1Mu0b8x+LuiElwEB3pVZZ3MSTYL
zrNBks+nq1vf5HIjYSQD4zZRNzT//8ibdD2x7hSfYTb1VyRrB/LrwR0h2TJZ4ZMJOM9y5qUeLu9z
BXDR1tFTmXKBJA9xQFwHSQ6Wa/WGt9E/mR76H25kiALyZxiUZpJc0uDaSHqUGz6R8ZM3SykjpS/h
HO1B7d0BOBaeejGbGkVvvIaxyvx4M/xzQQxPhkAwCiFwxt/NuDVtSa94mi3ir8wOgr32xFD5aSS1
zu5I1HJryKu24PTiQuH9WPPTxmV7j741nm7PNzCo5CP9ppna6j3tySQsmtu04cVHzp2+MevSIGfv
YK0GUzg4pcx6VzP/nbM9E4efu5Sgozhley6RnY833zIts8GcEf5bKyRlvb/dg49k0ccvYmS8mwlP
sfyy8MXE/PKgJKJsRcUUHbqWvuFmCsNXOH24pYt6xwrVrM7kaj9J+E8ILVec2b46MlaujiDHJv0o
qkO1CMCT4GGE/ctrCI0GhuWdzr3e/ABIlmU+jvu3Hx4LPHS7HOiUe9wsqbEJD+kvrKBwxEVtioxf
zMVJIuLWQfRdbHdNmUvCoISCMisIW/D5BbFr1brQvEwczIssZX1TGGfqfWipLvgEaTNDV/o/fSua
+H7CrH+HYuZD5+N1a6mJufsAY5l/EH33JaHQC8oW7Do97r5wUBPH6NSwl8b3fUZDkSpnpCPBC9rO
QAkM/Ouj7eTxhU+YU6XzfIyhiaCXHQ5NKIqzH8OPmReUQ9n8lw4O5sLWFi2VuBkmDPplLduME3+A
DaBs3bDWG+VMIs2sg1S+B6DTzgnNNUm0oyz6yQ5M05RfdKNDZ3tiEiOONUW4YkJ/bzIMdgbNCl2z
FB+XCtWH1oCfgo7aee6kS+wh0fsQ4epu6gRk+6BpWxN1bQQH0lC/kUHmvDQb3H4RdiCP+3opRDoT
QLTTzJltSrgI5z6T5blcq9TAQfqzqujgr3ss3+BKV1+php3+e4l8Dbv+V32GvOPYZvTygleRqfMG
PbljjJeLN9jZFCFktcfRhoTwtaQ+4oxqO8huuSZXIyT0iiqChAyQeyAQTSVO9d0+WqwN3GTw3YJz
BgP1qH2nUCeBNLsrGQgvp9vDbLNIu2Lj38ZTOIOrP7mD2NHtc40NJJgozwmMcQKptqX/UDuvPzIX
iORIF8tCaj3dW7aVHQsHweo73LoXfBF4TtKPLkwsYEdjvlISagcNBhm71Rjb4fQlT+fOxjpvCuEk
p8a7LZfwqmhD/3lT5AGAqxEXyMVAt1R1EL86PBlljCS/QnWOc4W97u751WRNLSQ611Kt2yxgzhUd
pqtpdksJVp4kO/fZMsyiESidN2bqZ65Ao4YRJmYUpyPoEbW0oBW3IdXhD0ZiXqqzDn1oUpFmoHfI
gQuPuCg1SuIznCrfYOVnN8b54GGEImV2alKpB9AUkMh9Xa/Ro1aHKHPVMwPYDibWRsxAy/KIAhdO
bd6lxRDOwTlMouY5r+AisxjLM5I9EBG13EhLJNsK9HoLwCTMZ8fMZ1PrZy5IATLJgAUtUVmw16lM
ranxGFuLLicsHZDjUG6vIZKfgjWUl4sIDvneE+iTy5hj/vW/XotzCqEdqQzV1meluXhY/peCNvoD
yeSYnuvRjNYhGgDlfWvVBeXkN04inytz1O5by/YbNVH9zc+1g9Y8MjTWV+wIGwsT+ec/9tpxkfXI
vmqBQoBOTK/Py+5JqGbU0DvdZB6UEJ7MxX6I+MCIacsomhGJnoNoocQ5+6jX04G/9GGLgzguARq2
5C8t77PWZnfGm6p78k1oxPGp+rPyKbdt2kMno/Eu3TylUL6OYGfYZhZsbuNUSwiDgvptidcV6u9a
UtQBnTTqAPO6Ekb/wrUb6ZWGCOIxp3RQfflFD5SYtwVYHFgOIqSvOziQHE5il9RM0Wq20zRbUUpX
TJkMtObbhSeLqLPWQgaKRQGlV/yMynOVF64XRZa8Vmz/wkuhxaQ6degB3Wiw4uWuY75n6VZOEQv9
jBKk9PQihMvF7OGQ+7BxbUDp+HmX/EXtUGBKStaKmxXRPAtuseA1CNedBMXG5uM+uvPQAhegpwaG
6ne0NjZ1jks7/3NnGHc4d7ErcVSfhjIL52MSsL5WldihiIUJCSezDhnKEyWeaSmCrAwMVrkKLtR/
wx7vJio3Sgk6grYt2JvjqX/1oR2b7FQc9n8CsG2hbgKafnsj8GHTbQegsJF1obaofqAUEhr6JGCn
tVxN9hNvhe6cSX5w7cQyOl5Sw+7BGMsYAjSdRtTGfWXP/HrD42Te2Floq1gXfCwIXaLTDLy3cL9i
3BTpmr7H0xfuxeGwDYjngoku+L+2xMM78zfhjhdpwzh8UVHZ2OaTEbAOnHGn5o0Fxhhx9s0lUnfH
/n7VGxNyXHkQC7L2SJCU7/8WysfTszZ9PYJI+atPt1r32D5Y2E4cfQzC+VUwHXbPdxtn/1woGpxL
EMk9HBc/cGZAMSwkjRflapoVmYPG4X+oqQKcYpYtjuUvphj/U60yu2/haP+r30KTDxGMQKRN/KTL
GaYBLVYebOF0ijaMfG3YL12LxdW/XTOFi6K0dCXEtcZT86o7YE+wc3fSEAT4OcjBxvjLQzSqOjkv
AKTzoNW4JsNCIOnQ4zRBic6UjOymCVwYrh2f3obK+X140iqZlz11OVpfUUBr5wDWm2hrGDT7BZu1
gwsaPkVY3yh04x7PLaUA0dMIuzxx1kliswl//jTqlQNxG7flE0ZyTeiIdy+JcowVR46aVy4Gfmzm
Tw+F0IPiBAKOZF4Msymff2nu7RaLJ35K48ce7/pnIbPaFqUhDIuDw3l0n6EiUj1Bve3MUhJXvATo
CQTTlP3vfokad52QVQMu9eS27oue+4RP18fEIsmckSpt/LytKX2aZeGv9hfmN7lXF576lF/+zWeC
HORmcdxdCQC6X9pv4vdltcvbi4qg2Jr9U9go0iet2Tyq23+oFFhiygmt50QlzL2WBdfOVKUr2DDk
n9OeGfP8qagclN//OaMRtbAxzpdEDZnz/hRldlJCHKievvezLlE+Iv2DjhwZG2l5uGb2yMBt4wEW
Gryz+1DsMfCZF4bp5G0cy91PDElit1zYp0/W+UEptR6tjNlyM+/08xkZPwjytCmF+wQvvQEGxoZh
uYJPPWAR/CIgvhatcCe63owF9BRB97J7sgGIfJBbNwdhM4yuUQXYouNukA2Ix0QhMZ8tVZlgL1tj
84npfkhZiNzIuWpNAQpNmBCq2XHbsX6paeCT+5ybSVdz60NUuXZzOi4HY2eVkP0cqGrpbY+2vnBs
0s9wYnJzL7GNkV4HsoCn0nzImDnSYuYb+8/xiK9VLyjsJekA8pVmZrqezbiVaorfslrxqrLsVpsv
Z1RoKu6xjhnDLVqQ8zb7/PjMQ0I8Ks5hzIeqBmkH5ll/J3OhW3EMnZVaY7VGvK0h4DzTyxkwhmRc
yGZ8S+ABYIj4nkWsJHCEExwo+AdC9e1wisGC7CI0hw6kAt+EMvq6FAHneBcMMswPxg2aGntMX1ak
QNJH/lxBwyP5SXIdl0dQnnHLbjuEIe5g/0ZZhAXb9lFDXoi+yIDzzdAAs6lcvABrCBodY71l1djN
fYIRDHoMT1COy1RR2MWxnaaw+U5iTqjobVQbExbjK5PWfHRtRM8XlB2RO12qOKA/d1GWDwEfH8Z2
LKfDydJ2NbAXr3FtyWC8cicyhj/UOd1+wsMRpOmArIA6+iHjujJ0McajKUHxiWJw9m43GzZNedWa
gvztl7owyAv0sxOCYfyUEI9LixMysJcH06i+/EyLTUzfqgm1wifVbTyWtxWxR1yVO8r4fZe5n5PV
FTua3Vsloo2AaprGzjnt16mpGO8VqrUkM9TlA3XB1i0W+I7Djwk+oT+nZSQER5lAqQCVdYco49A0
g7nPICdPc5FNyxjNug9v56jsVkS+jo6wbTAN+m3T5jeOJHmz0wfEETbGmOkDp6IJKvyJPxy/eSz+
pDUR3q0v/UM7udUV1Ciuki86sBKRCXt/oguUOV6VANX68U7HE0kgaN4ISL4TYs7pKz5y59AL4naQ
0GcTPF7h8ovGFiwZUuVs/FXGYWL8JzDlhKpLpUQ9BGZGWItyZaOtECU3oJpwrcrIuGfBHCjia8Uw
+CjU97Fp6srA+wjmlt/zFHsf2+/bv251B7/SDwX4zz8faTrPiCnh72FImC7BB1cbxkG3ku4d29i9
CCKl9YE8h/WU39RsaqupRgaTcWSjVII2UouEQPPMj24Js9zmMNgdL7cRX8m8twVjolzkJd0b72Ub
g5NVNzH27V7CAeNtKiIBn/m5VNpEoh00Ts9cDhtJkWfJ3+9gCj1SAy3Bh4RcgwE/C6DJ7FyIIhpd
CaxHk1uRyUVPqYcWQSX2QnTAIxBlqBmYOuBpMAG7L5C7+Kz6KQH1Q+l6dKyQDIHAvywhIAfdnct2
knO33OD03Xa2Y2zDpj1/7CePj0xfC3Gbcuswpt6VFAEjvQIJ8Wb4xf3O7UjZyRuw5oJi/0zg8QuV
PBoHICOgqUB8o7IIoHpTEfpAW2Wx936zdRHOPCthI2F2hMFk50tSgYpqkXB2zGqWe6qG0BqsVJU2
g1oVVqmZUdt3dw15W5bcrWPMad9yU3gDoFBZrZuIx3f52z+/bSGs3gVC4GV7Y2DdKz+LiGy0t7cT
9+gtE3Q216MQ6bP+8uR9UPTrA1WHYJFpkm2a1c63qeemRWy9tWVfmHtqpIixryG637qz/Kyw/jEr
3RFN27UVm9toZGmHqgDGK6Bq9mWKk4tUpY9+DSt/ih4HLrsEoqBcO3wAss0cFhurVaxERawVeV8K
N+scl+F5m6cqeWix0BeUi7mb5F9QdQavoaxGHLWqVZfMysaHdw4JoS4UMLgH5ri5yVkBrjVAOyvd
j5046rT+QSoWXl0Y3Ms89cPdB+lDIhoacu4ELekw7nbAXlzLsWrN5Rx+sJ5FnBdlf6EJX4CzdnEW
g/oGcQm1+k6/9CG7XNuj8+h9aiFkx7bJG9U707EZRQkjksaw4jgQJYGZ5tO/F4ecU3GIjOsyd4Np
l4jv1nKh6rFWR9nc7ZGaLr2BPUcLoApgszaXeiVHyoeD7oEavLsImt5vQuO8d0m9G9LQuTY2wobY
ltQ+oaMPOAJUUoLmVzHyO75cypuujZm6HuC6ZdewA64tFjWK3DnYHal8WoCvigJvIFNw7GpPBxYA
nBjOTlyvglEGTGfJjwUj9LrHiVPg89819mN1FmVyzB6e4Li6qW3usqz5uQRNFAJ9KsYw1AGtukLs
feLEfDzra+uglOUZsPR4EYjosawe6FuAprKMpudIEmdxiRD4EYCgCiplwh7OvyVt+5bY5ganTTPR
t+GWXhtr2czy0H8jp/YxcjooNCtTHPUJW7nBxIktrWbDiCc6xFnrWGElRtpyHZVecxROj4HPO0H/
LmRs9n0d/fvj7JIYbEYOlC3yinxBkzStD5f6URrXWLQo+t+JSHGPvru+Nvzd8TslfXMnQohb/NPI
gnv1G+b4sWZWl24aMJGB0nzbNdGBfPwAxWoE6UA5NZQjGseTVPzQWvaxMfxAtlLSb0ghugRW4cvx
FSnL5sE37eBZpXr1tCzZ62O87qTIR6u7R9ScxlgGCkzA3rYmUwCtssh4K405zDWMJFMJlM0mvlHw
gyc0zW6P2HmWbEu6oemfBC8TnYEHZ3n/EsYihOssUkJhEBsMQw2NVCIXfIe5EtQeX+6QImIZhkHW
jvBZNjvSdRRZUrLDXsu3xhX5ORXZbsfcE/4GPjFBBrf1lU1aAZDhkvM39Yq52Va9a09LaTTv+kiT
im1Xp1ZAg2rfoGuCefyVSarkpamIv8xZlin0idTF6p6JPAmiI2uB5xIu9cdisL+LpkILOYJjxTsh
7psO4fYFbpl0aGRFPVMP3p6L79AFDwsNvkZ7Lan81hy6EMeK9Q5UfZ6xRWNyR6lGAqAQsmugckXW
bg77hv2/1SmqWm+VAM6tT2FsIweO3WZEZVCISyFcQs/1nLhZalQXmTX4htkTrHRf1duZdB2nU4d5
wTv63+wMkiMZVnulnovxB8kynw1NH4pwfeUeeAFfMnzI6kBrw3qNJ6gTf+mrQsgmLsMnntsC1o1j
zdsvLTs4Zx6sQcPsvhmq8nXZDC6anQrqXrpBEv9ZHgNpWsabTZtGFlY2qRBVSgyVPohawn2OZh0Q
SAcAHZKx4o86wcd0EYBYQLofEUqXg7ri/dyi45coBFe7q6Q6Yd9uk+0wahNK3ecg07A3/A6Q8YYF
Mu4w3auYr4v/rz85V38VFG2ompByrUKmVuNaHdNb3TWUkN4zcAvrEJ8fkZN8Szu3ITG9V22i/Vl5
JDSMP5FirQVSijH0bvBu0QtQqc1kn2QLOTPM9q6eGAr/SqwhZRHKGHl4AemCn8EXLFFMDHyJwFuj
NDMl7p7x4oROD3I+yod+yKhoPU2OUq3SBBBAwxK1+hTFwxuhiuPSwVGw3qR7vkuiZwvxRjRIuhky
lqNxtAqxROdEeMqPdK8SAvxy3iQ5VtRZ+p5EUjXRSe1u1fqRnmYY9KMgJm3Zh00IVD+w+60Zspob
3VHVSl1rZRbVPGfRBXHCpl0sYKvAbid1+8DjO65UaX7Q7N4AXqCjS+FWlPuhbec74nw4QBvFO8iF
yky0mq+ky3AIx1UHQHNztMK6p3lVkqmySahzejsg3Da2YF0vZzeJc4fwA6hfHFQFcMY5NVjcoC3d
F0sINxUaak2uvrUTF2nxs/fw3Bere1i0aVeH0ggrkpC4Y/ScDNiNKGLjNWAYPsh46BjAYZX8zcE8
4/I86wJMhwMSpQ5+CMiPUJ74EP0mXgQtvcglkggVSCxwwMS0GkbCEuOA95xEVok7/9Gq7s0JE9vX
eevJR5spQY5o1eKeSAdUgEcZ+SRnfm0FQyRdf5y6vmE7y+uOBWyrdGt/Driy8jgGUWrsTthyfb4U
e08LX+Wq0E68uzrL3KHzYA5Pt+EdzXWZe0mFR5bkUIYCEBBZRnkY9zZZ2Al95YYnav37SNByC7iK
XP7h2Q3U05sPMEqwQNjsoCpOKqFqavsk6ORm0AysN6ZY4jUS935u/xktFToq66gZ6eVCvYqhcXTr
FHbzLyi5rrsI6RiHj0DyFYVw09LHs++C7agNS8VYmm9WegY8Mb2tI3r/t0JojTXgkxH7ifaJU/8T
eOhVBcmWLbC3x4S9tQU1zXDZpz7bigv+QuAqaOvVtC1l407+nozrILQ//lkHr0G4x909y7o2CZty
XC1DAaoEosdad6TjkRt6da6WUZYeF+HWB/bCC5eiVic2oiLpRe/DHbJOOP20D6ic+7z9aAKShEwd
06A2fJxvYKc1jDxLHUil0RedBwKcQM3kTtDdKBW3iWzNtd107EDQBAsz6D9K2ScgWLfWNSm9xybg
56pinS8XSQ2gWrf6aNTCKXW8LmT6abg2VTEqIeS+d+17pJeyaMvkEX2hs/s8CvhfCJWwQB67rA5/
8U4pfbeNN2Sw382h6O1R6NsfFUWZ+krRk1iLvg3GpvhVHC7vrRdz++orU3k4MBFf0OOx5LTp/9wT
pfyUnVF8fbaNKSm01sac0fCAlKn7tNjvD6CWhqZ14m++kag/Nk5jiiZPatakpNfC7wblnAitO6Qf
K7hUk4Exp788Qrz48D6dzoY7/f9+YQHdFsQIwmeIAMReSEizPajiHoRvTo7Z59kHKJO6Ib/dB3ZN
1mKYi87P62Kvdnj3RP6pm6YAzwXeFlofkpvso4YP84YhZp8MDsJCkmdPqE2o4vYSm6QipLWe4zqd
1qR0b2mD5A8xTEwbnOuUdxcSJ5IHBdUypASkE+eXNKYp+/APiRoLeZ5tsGifh1QU25gafUydm81r
IVLnoq355Zsd3lg9r+IUE4XGaWqqRn+RSSjwZMqvnEA6Cx4pFurA614zK5GAKAapLLCmX7ZvCSqT
IiV09zgQtN7K6WDm34fvPlfj2nAQThq2q2iplHaM6yAgwzs8T+hRlxkaCrtt8MqPFIFtw6UJRzqK
rQDCzEk1lnWvzxjmXAlimG8ijkIJLW3joxejBKEfH2bQa98RidSjYGma3J7O8uE59stp/3D/HKBe
h4NvjyCcjup8nfskHUj5SBMQDsmvANiy5VTJ4zLz0WZl1Vwto8bEPtM6bi1Dro9UsjEk/R+/DZwP
09XWle5xtmZ4e7wSpVNTbMYYi8etPqWqC+O1WNwXjjXx1Kx8VvQBRXMO50m/yg87HfRjtAyxgkMC
Wa1YcQW4tJqGux9Af52U9eBmsySbKQdNxDSDYZPmAGtWAnwnz28AHb3n18gVv7EoxSkap1bNE7+C
lgMcaBoPYxUmwdjhh183TyrfMjuHKFselWnR7Oi/MU4N4093ksckbXvk7OaarRuzpU/vVeef1xCa
xuV56G2M7PyKKSsYQCjktujvvff1gt8o0tOsvLtePEdATkMkeXQoZvQL/zvC/g39eEKsvfYbYQEH
Se2YSpzxnAM/piXmyOZQbHHBfEuf3/bOsbtn9UwV2Lr3zE9z8HfxRrTNjszeEJxFklSLJB10SBmD
Jx9xwi6+N7s5/0p7F8/6g6ZYN/HKpxHyQ2UW4vygPNCr8RwlTM9ILmD87/Mz/aoNU8PppAMFOnwz
T5XS4i97bY+27KfzSCF61DxwVyns1jvCaUEF3++iEVu2+LsowJxDR9RA0aKrFDOvZxSlq0pnzDS3
cM7x/NoBOszdf1uvLUcxDC4UuZFscVdpO0FvV+c5wFUeUQqmW0NYGn8WBIE11sgG+5S9C/0Zvtgy
GQC+Ew0U1IHDDe6ZDiCs48uhC2DduCyMy1qyAiBUi39UX2NnMhfPfr04IK3zt0J2x2DIFbA/oG+4
SRxNjeHMCeE6uco5gzJjqm1/qC1+9e8QUNiiTDxjKqrlXusbt9xrBd/ficcLNbElOPnTv5wx+Oid
QtH1QWc/U0ZUrz1CQyWR2wUcRrR43AGo0Ltzqgjz5W9JDwqMqdkKuRai5Jwydeyw7LpjSlpFQzRv
ZUKMHev3JN+Pkj1C7SgFImfNHUKhg4EV38DS3W1YKPYoFZKbllaHs/x7L5kAZonRq3POSzMvfmCd
j7o3ly8YRmIlJxNFqYILFHIEB1b/1KNHeO99TmG5XftQ30Z723o994PfYuv9XsPc+EvR4quUz6zi
RCzrF0Z9yexk73Ovfulr9/+dJBq9OHLLMyjqAZAoZ78rqG6rKvqNmCSwPzG7T7zWBCrucbgbYgW+
NxdpbL9L8P8Vr1NITgWWWS5UKOktv4lDtsCJvAYUgy2NP06KZrB4yrJ7lyi+2M3mjLpD3jCUYphv
/iKjwkDFCmrXj+wE+MVjKcksZI/VToopZkSTFGyJMODwrDSzmzUNN5FQWM1gtjDpqduSaTTA+RBk
Tqo7flb3uuBeyuvcjLDynZVGOR9wZFKUevwOPWZ1VdI2MCk9ZMrSUHFCWL/mWf/o6OmlUEK71rp0
pHoeE6FUt2LGC83onop3NQs/xZTj9W2vIhe8i961Hc9nqk94GWsPtLenDSrKBL1pcSOStJ8HVbpF
CVOjOWhaleejgndM2tNNU/aNF7a+tTsVKkGdqp8irsrd/+V8wjGR+xvO/jOFS/itTj7AgIsvqo9q
HhraLPMeUGpjK7YMkPXAxCj17doW1K1o3aal67mRpI97gV5qX/yhA+SmkyMo88oPtbz/W9VfbcC9
4/Sv0S35Sszpx6UxX59BELzkj7pnYCBhUMu8nez0wksuNVI6YRauR/VpBlIcrt/3UwJymegvTyFB
QMGdtVqOHsXffL3CrfwMQgVdGfw9HUDXvh8FgCYFGuEeu18tkIvTbar67g+bjuzX0ijhH64K0Piy
TtlvewDB9LcuER8g89NQblS3/V99W2Wmhsh7ICEWT3ZtT6t/H44GOI26TLHRgTsRYVkLdoBsBA0w
hBoJFu+tnKP8YMowZK1/w2EN+mYiIz7bSdltfutn7oWjhCjo0bwQJTDcrs79j9m2nbfNuvhqL8kv
wrsbcN+G1EACDc46YJ1FfuME78LSKL7JuhFO/XiUz510sE0qHT4cz8yxkVzNH1knKije4LB4ahhM
SWdEM8CfX8dZEkVPX21M5EAJJY+qx2fYCPlqac/J31IJ2hkzn+C/dXmjajqTcP52j4tfUCTelsxV
OMX0Mpn/+UvkEQUnhnK/+Y/+tRHnAz/Z5YzGKrTdzSQvDcxYCCcLIoKV8zmBlOjCHNFNuzjDuQdT
J66rQi6RtvBEcL0sc5ZeR3PB5jcDLiVKpxrW8IOBaFF1+13ECf9sWDxn9lzIi8uzqpA+03lARtR+
ShLx0FuHQO2GxRVDwD6db31CbIV+SVe0u9gus0trDnmUWxuphc6Rm3TYelE6E3XRzBaRXH94Pff/
y8vJt3SRYH+XeR7fcfo0FB4I8lLmIIgYc4zGU8tL589iWTAU8DSVeJ01X7telkssZH1rJcCfbCzA
5EHkI1VZET8duQLBc7HRoNbHeAqjmYLefQb6iGxByVnf1dbOnaeOCMz8NNSKZLF056+22XNFYdEg
TfyCwc/RZ/HSzUML71VvXLnLsz8PZ/MWVharo9u73QchX8NnTUnJensIgvNJxr9TaO2qzoCCqcLA
PKkUSjeCKHty2NFmqMMpBEn3+2x9ves0ryN/6MpP3jezehpfbUxVqKBlcC2VEEtenC8F9KykWYGi
DVIaIAar++WiC0jJQDX5dNBQOhXdGqxOAAWWj6x6sPvsiKYRGmkgBSAgeRHk8+Cjxm4Qb5V2Bd5M
hrI4ufLET7CbNu5pZDLBE8vS4KAZ398H1mY1Ae0qjXl3qEkd2q6Qfceodnz18DomLgEVM7pIS7qE
ewCIFMvaQ8qzIdq4X+yxtOvUPC7pt0UUi5ucsJgVeNPg0yesf0EzHhk4gNQR3QPTpFnT2dRu+CLc
hbPTqmWxQ/Buz1OVnj4YHKCS8PcRS1w95bcfvgY6ShzDiSAlId+0I8i3JaLThEkhSaXEocd7Wx+4
Felvi60ZLWMcwwIG4xb4+ToZ8DR5YJqT9u30QykfNco9Pqhgb2HIoo7nYR6M0UXglPbxAiNjNiXr
eIN+liJ1xYWDyyC7jF7BiEOzaXqCEtjgPp1ntMxwxdptnvlQ94yuGaf2oMjGA5waUmiKOHJHE8jb
zz7l34158EKWWNBRgXA1fPlmGEEfPzEA/9JA5FsdXZLvgJdYZ+hVUHX/gIZPJLhpbpy3E1W8/4h8
o5dRmhME4YQ5XmRwwliIeGdheJwX/5wtWmSWoZBTcjKqtAQnSgPSEZrmphOJXLGogB/412ZwzqIt
jKqRpp6V78Ph9Xd//A9QT+dYaA5mAe8u6SrDWski3zAbnHqfQKWyzlkERT1ugWbi6X2TNgDrUjKU
N5ODJwzjOQ1wqajJOrUMnHxsukWm77YH+/xq1eW22YUMrZ1kF8FyPapLaHaDwvCjsg9ReX8iFM2J
eSYu38nU35TejQFUlGVwCz7K1jcg0wndfz/OjW10RbSWVjKF/bef/HVTOHc30hx4V3oK0wrbNm/N
mKY/MAGkYy93h5HoKbELQSjE/8ZE76V/HKWtmFI/6mrchqHF4jAh5i22DLWzewyTgPbmcb5kQuW4
/I8HdNhZsiecXJu9q+iUhYEzwIYeISiUqhgi+XwisYRMSE0NQZGCCOMJVOlXVgmJU1DTd714NvoC
4GH6Em7wcgRV54HkKdQ6lqhFwYiABioQdWgtgJkw2CU8uzhN0MrExNyUoYV6REu/XkqTpvNQ7j02
z2jN5pUk4cvB8TxproYyG8GNJ4OilgurEPq4arWKPDKrEK9YmTGGTp5Ybi7lqVHKgG5FU08Y4kQW
rt3nahN8xpF5B0uaryQfsY6mKWEBrkJ2htPTpeymvbXqBGQ49kwp23tN8M4+oqXB3NotGpF9kziB
tfl32iKqo9t3Ts4F/5i+v/N9SGhja4a5/Q+vdvvQXvkCtJ0+i+IirfaIqVl5yEn8red+uRDZ1EqV
EW11KlX6DmMdpHAiF0/Sg0NvSewi0AxxQ9zb+tGPHWhKVExeMyUif1lq30JlxFAzDjcp68Z0u8EB
KIfFZLNiCzRH4cUucJSYKcBQoIpZ6mwkYUspvOAmIb9mixSHaKVmM2x9QyRjeZ5FGE6BFF5gkZm9
RxeR1SjsbAvGSc8uyIMUcELbt/6rbAdeSMDYxXI6Bj0zaH5NgMrsKKm3uPKhjGLMXCDxiHj1UAZj
wt8BFubJ3+UaPt/kmjOiIMxGNRLJZKVrP4h5Oi4ll7TWvKXqDbooqGCwmQeKYEOVMS6PxTVr9Hyw
uD6FZmyt9WlADdtCTQCKVlsq7QtDer5CTLV1CZr2djNZS3G8O6giGaDNchFqiEI0QMGqXvAdmnwJ
xcBJuvdNuEGQWZN7RsEdABii7GDCy57JVne0YW9FKE2dlWdfx9NA8MCdAR3544PzfmqMZlt/prLu
qmjpQQON9La/YuhYmwFeDTL2at34RzFj6mD/cHDE4yLratMZyGJ7sbveXfbzk3vorTFPni/8TQvP
x1OGBg6qf3lrakwITb5zWFFeH1j1x43Eonum99TcndsaBpdvoOcVN6LaFf7TK9Qx7utAIVOEndMa
qpOPbyc1b/xkffPZCFQqw4BU8+rlgLOu6yUwRjDgBVzgWqgVS63Fu+vK0KTWaavpCGUgYOVifmpF
vOpeIiumQ7shtfQUMMB/eSd53wcxp7f042J1Gp8AmPiCHc+NAs0b84njpTOliO9AuP0S1CE4QYXB
9SjKcN6FnV9UgvIryRMgMAkkFl63C32ZNisL9EkFnUegrmDokrGa/UrSkDChzBKTt9vh2Cp7x5Iw
Pncd6mSplIuZ1HXMgKRxjG6g/g6NHYkOaoJB8tawiQu+HpZ9gQhIBzAtW15FqOqijPksg6EB7+yt
ytUflRKyN3LE82iq7mOP2ggk8EKjgibd2zu/jhVWCHBr31PtRNz+2+EHvZ2Gq5vMhVfLXVZugU8R
qRdlKQXheBYzE4hJj7mqSHF7n2RVG5IvpC6V/oyXoKulL2Kh3VUJbi2fJRIS44fpo7bcj0MVNs5v
CJOk74D2h9jPZjjQi1Di8KlXIK54rlHsrzK32m/1Deqc8PqRcrMcK/G4cL++FYMA7m28jqg1CRKt
pi628VshKmfJFuBKpTNOBzzx1otLD+0w5HJEwBoJeN2srsR1Bm0hBWEsgNgM4PQ/uTYnpxwG4NXv
crJ+oRD+pO9GdE4xxJGSC96Go7OTJ2VB3Ceq8S+bRIUTP0r23GnnvqDk9olfxFnncssMBT9LhwRQ
37+aLsLzhZT6XIFPxRQ7AaACPj/fIHgwDSI5KPcTOyEGTS4nV+V24gZC1CaNVFcdcZoUWTk4DLeW
dFWODRtbTv8Q68wZ3vQEj3s7DDxA6t21nVbZNHTpwpvpcUx4JdFXOzEiNuGQV0ZbphOnhlPfiOku
CPc/M63NFENI+pwqfXqODz1rdx7E7OqFcOIlgqPsP3gDDeKizzjt9SJspm9p1k2wdL7NpgfP1g7/
u5e85UO6Jz9OqH3IPHlN8O0t8SerpkUfX4afNXpdEyM9RpWb3zfgulp/8f+/3r/TybLOdWdf08wn
PDsQLT3cqW/9rvbFSDmcW1UbHdrGTXs/19aE3vLOfxo5Uj7XLD35pYSF9bZ4MUIJB9QdEu7P87pA
uqxeCjM488ckOQv6MQnRtvSyIiBfKQFc75m5x3H85hrfcHz3DBxw9m2SFtDJ+ollj1PLZeq838Qe
xLb1OvUPfyH/mdPntJm4KPo+6m3yYbhbj3Ho9bMjlsr7wXbPqcHfep2j88hEZn+rm6k9G2PKez6r
nM9BphbgtAetMQYt0TrrFtbuzh4a4S197izq4O+2tK+64nSBWqLR+WuYh7JHE6aH85JIoBt/T+54
tjZy9saqtdH6NwGOftSqhFd2IL5gTu9jDLEcxOhAV7FDyBcnvFzYyjocbY0tQz3McuJz6fXvOqPc
u3ZrWA7xkvufHxwITuJv5b6t0RZvVQyI8yRkVWvq9wjHwQ1pA5pJa8M68NdFh2flReLs8mwq5qdz
nhzFCjkEBNDIJWyQw53eJpFtaDUVV2HmDM6IUhw0oN9ngcpxXrHilSuDlVrArU3st1PRK05ttbGo
zAMyNi9j0V+XhNvfJPsD33RJNuReroCoaPQKv0eA5maRBjaj3WpW8Iwzy1hmJjo/4CGTuaBbRTNr
N/AjaiThfMQupCyQcSnnK3oTrn5QqgFJ7WMvfChMLkKLePYA4DORKkW9eKJkzmo169z9j4u7mWUI
lnCRYRSjUDcoRaCijoHsBZcuZfHS0OjzHqbM7gO3GDkyGHgtj9/8alPquSea4QfJfCDUjyO3XHQ2
Gn0UA9qrUtVHtDIquyBWnotWJ1NeU09dYJ86tZL0lTv+neRI55UtIW3OZyMoFoxKYFqyA7pcWJxe
+y9ysw+hQxVh/VjshNqsxPjHHy0psQFtvvDY0u1Xo34E2ftT6NTHv9aMGlj7ZVvrntgoKMHVhQEF
jRMCLRjsrQuq2CPwKoOwE9PHYVmwHZUiWpfsFNVqQulde20J+oM/L2LoZLmctAmX8HET9cCy7etX
OxRwhUf277xw3vFKT5xlxsGkupZC6EtLdG3JEKSekINYsNAiFXDoOBMzxq5S5XZ3jVWNqQAAkJcB
1WNhElQ9r1HYyWR9xVWKa/SxSVUMcWN345mAFqPIX7eUtM9xNAayfXe2SpIv7z6LghWcSbkwhebW
B4cKkdHh+1zijXicMpSQsYoc7Sh7VlQqbnNVDmOhkU0+eHDmvYLgxMK5Fy6vkyB9+aF13QlfJsxN
Pn0y2h/NLXhEUatTHELAvSIcWIQ7Ugr+rw47BNrJYIoVCx0Gyr1wi97fe6XIE6YbA+pB6B+QWJ8P
lyUhWMkHj3ium3I6yavEpaqvW+u3Lymyft4eHrxJ++UBqoSBRhcV3YoJdRyrurv4MVzsF24iq5nw
CFG7f41DUJ6vZgMeIdA5HlZnzA/1sz025DiqAoRI59pgYF/wmtDzZ36JPR9Rd5XaAj4SoQ5JNexd
fN/HwAQpWbSw6x/IIEB5lCEvHHixnPPZIqRCUEJRzhybw1I2nN23rNzKoNmEmJIwuxhgCSLuvU4s
vrHEtiKcIptGnYhIX8r8FSp1yPx+T37GqBNXTlzEOzDBdOfBVgePlAseed1hfDaJXZkBnWWdNVmT
hNnxuXmGheJqNY9AvYv2F/84XZzG6qf1I7SlR9+tAMoEViMw7pdvuXkOaPWqld914PSQ+SfzqkL+
8HjVEd2yL5RGyFGc8idJEBDW+aF8RVbvSywrki7cEOhZOqie0eLYsp0fnMTSGzcLqfHppcUWDKJI
unPS4UtL1DZxThXbcPdcPR1kBo5ahnJQZdZlzfzllB2WcsLEZYootngYBiH5Cm27FOfUq6gdHT7w
PAQ53UbgxyOAvcqQJBdKELCKKJuuFaptuJl+0RuLE6NN/KEC9leozgIBBRBoOE/r3zsOj31gOnwI
Z5pwMznEi/AyVPJC+AgzhIjFcoN2kdCvA6y01aoKPZl4VMYCSy0NHVfLCY6VNkJJdTcPnOBFOOM2
gyfTjOPRMQRDIBKDWOrffOHBxH/01fKABX5aeIN/TO63Ru15fxK1NTk6OfckTY6+0no5mshcZe0G
OCQxSsVf9mx3ZGR1Bdmo/GakZCoEBEVruNiB7bvpa4anwvY0JHPZYJhkfgzbOWQa40KJsXBHmDjO
N0KFCb/rOgrsXIBVr0rHUSUFh7jQmkM+8f3TV/TtwMJ8o/PaLtcs8sT4nIOSM/0mKcaT5WUXtnoY
3Qn2hyv7Z2HnZDu6o/Iykf1UArEsC2VVcz5qG9jPOaH6jqmpYO8yZ6is5+sAQASrPLWA5hGd4NmH
Q71gaVVuNi81YqDPPjeVjaUmMEjE68bzYz4SA96mG8IoLCSt1oBxK1t+unYza/fgb2DHHBDjtvwe
6GTP77FQZ68GdhUWhyvLIvX7WcH/nPRMTsDio8J/wSNnSXSJG1cUfS8vD9wnQD6BKo92QM9k5JY0
vKfVzdW2nUI4Gwq07g1vhTOhHMBtWWp9GKRlQYPgvuOQd3ldEM9nW42KXgcY/dyQCAiHURVaOqxN
ysxQG/MAyo+uE4mDhLVCfoHrjeJYUqkNXHaBqM+LGJ1QE8/9tAsY8tKLxoMJzJTZw2j45qqYXa7Y
rgqQYw1G0PaoXrkVxPeShJnSuK/4HSfpJ7U4HpeIHTt5oedu/XvTQ5+rBxqogQoepzmQF0T0XNwh
p2HDV2q2uSsvcF0GzZvToqnybBNm4Vq2AtrJPfWmNt+KQiLiJ4s2idal1Xq+za3oJQbTvjhWw8JA
VR4qrgbjvSqSjMytyB1EES4xPZwrewG+E7oarBqe3351n3xBV61iNJ3Qf0Itu/+CdnY8uhBMec5v
BoJYdAcemzvOveAynx1F2oL3iKRwJ5nOMMfvHatIkZvB48b+gTo/f6WFRAmfBb58RK78KmfcZr+e
8ig+xc/3nqXujhhICWoz3yX1BVxlUwLgncfIeHujtKLnEnRG3iAsVAThCmaEFmURYiQiFHwUvBvk
zLgiLpxh2wbv4gV1I/vlWeS5R8+qeVnNGNNQ7JLcNl/gzQFtlHKT17msqseEcpSQA3RrffrMyx2v
0SMiw+GDGmals97QIvV79x4V8VGgDFQP7jTsnw+rb9xV80xDDxjnjbZRQKNAiHtQr+S/sYQOhzvz
Uaul6JAGGaRHGkPUmCQg3DeKJfwdACVhBklVjCeTTjSqtLRKdByEaRpV+OQ/dORQwyN96W/vKBhT
ZjyQD/WwV+8tLbKLKskOGgu8c9uL+rzyhep88XpnZyQ6BS16HShzwo8D5ed9kOkM+ZaFUP3HIt4Z
Io6oVewCsWiiX/nS3NPzP/hNNVPtzSV+xiYLVdFGCSQ7g+Z/Ia9a4iIgQpNu5Ak7VT0fmxYadoUg
YEuNxsMffQJqOsBl8JAYa+TL9N0dV4Grr+qOivH5gllDHila+vM+1q2A7ZXmW05JwYQdJGpW2Dgi
1cAnu30t3OcXuWIoGDSoYr/CYa3dTDH5YP4lbYrk3v6WVQcpyia46YW29CirT/yhHFHN26zdOvc4
XGYLlTPoXXbms8a0gCtZTx1l3qxkrS9YvrcO6JdjnwI8HX4OzsfD0VfflQmR7U+5D+Y7Mze+SXqe
l5yHjd+BJLWFHaDALElQhLw2fmSD9pdcs8IvS0deYc3W9pBni0q42dkcxKmFVqKrJcgbdoWKSnDE
KIApj5tNyRvwFjrodvHIpa73/pawlpOqvd0QAj6FJIGdffT6YfnQM+M+AwyMx0tFvlYagDz68O9F
OidK0wLuhj8cNKmAFfsPGHmWqns044zhwn4F3HVVmTS92Ux/Lx2ukIVR+VFOJssZW4ks0xDwwdo9
Lz5Dm7aeLbQ8n5KE6dl6QzkbKYLhEpoCJCXFBa1FnOrFbi5Hp2V0E1ux36luR2vTUmccH2aWUTA5
yqiW3nFXZ49N7/ryHtqpmDso+M2uvUatZZwMRl6LShGKAEVlIZaYvAPdOtYhEyByi3idKc8xVoV/
99tc+uYju05Mll5yGAjG55QD4gkaJ0CyrVUFnbPFrJVFMHp3dn4jfTtcAkG0grQpUaefznxVk0Jw
bOqMHIxzntcIylCXUkhj3eSdy3NKcKH6CDgeaXYUDmT+ziopPfV3vCKVze+CXR99FNTrBQkfj+dL
irSK2WU8xQb41N9lpzkM0wHj5AU1GTxfWHHlcojeyzgBYBCZIOLgTibtpSkIOnB+CAMypNYHq3PS
+FHBvRmgX2TP8ySIAuQTBwJMVat/KZ8J5yb/ZYMq6ok1KJJm/vLE4qIr60k+z+eor9jXl3UahNyK
MeMvqBGN3xlSUxLdBwsmNkaSC6w62vFz72mP9xAcb1LAVKbI1EIe/TwfwVrqrAIObqcqEySKw+qJ
PJqPudt8D1/KWLivaUxdUcimqpnBgW+hg00odCT/uZ8n7msvJrYp3a34DH788RRr7ZFfhoMq79Si
gf/2wg8YbA2AvKaTu/iiP8b8rApweB3GUW3ZMKuTM5G+XDDp8LADYkdSz1XwR/ihlwTSzN0Yo4Lm
kYTNu/5rkzxC7hIY68iymrgACiP8F3PypSXMJvxUURyj7PS9WPpr26SSi6jjrsTIQ/tKMVb8iIkD
u5CVtR+98dXaAPwKWpucZmlMJb87GsXI4vSdnrfjk648j7rBjB5ynQ6b0C602WtgavEXEnQnmaZB
QgCEO0uTpzFeO0hLfZMD8zqoqiZQHyoZ9g0X8W2/IJ/bhqfTI93KXlgxCsWOjvHzbLNta/9sxhHr
GEe3W7RtOjBTpznJ4xhfaJwqG7jdcPcNPt+h6ccQgabR/0Mi3KhYcbAZ6AI+OWpjEuM5jhM0dD9w
nogQORI6L/8qiidPDyy8QA9/Mcw/G+Sdu19ydJrAqdZ2Y3jphkANYsQfZw3ayFUunMRCThImf/Hc
iMAqhHjf4oW34ulAkX+yTjwmwuTIo5qvDVdEk1FxocW8N/yy2R8cCTHiDslgTUxFsBDBekiTOULY
8aU/huhpWWXhXPpU1WfsFCaMZYqkir/AE3vN8JHdt+h/QruGpmTdtUuR2vsd1EH3JrJ3H4fg3fOr
mZpdG6Tb5P0rGVRnyGIayIg6IAELRhDlOjzN6BMJAlqFVcv3ShRAHZDH+xn6xlT6f0iEU8B3bMP1
UH9jeHI3M1JsJH3BxEJ33glM3o94NzO6BlHccYvPabNR1XuG3aUbs/Suv8i2ZWdwB4VjBMoFHd8t
cx7uP/To4GYfons5I7ksV0Uu9+h62Bi0RG1Xmk1HHkuDs+lrCTyVCPfUZCulnV826N9zyvca5zUd
yMbsul8g1f1tTdrEOa2qWoSxrD1SNUXc3Qco2Fi7vEU7fSrBm5A1JZXWmKJrto9jM+d6Wok9n6EO
SYFaVErRYbho3/hSyUBKHj3QmQpUbmts4S7KB9yNYZBfl2tcYXnac01459h7+8NO1xLez1/2ZwjL
us/vaom4K+zRmoH8WFtFBHhZVpqRajGxXn42nfqz9mm8DuKUSJta5/LQQGrk4ChifXrYhj1rSs0o
Fqc9RI3T6oAOmSBhMBIN7FHYmC+/FpLmMc6/2pveOGzFvKbKhfXnjXCvOT2W27KABKzqmtuVZKxK
2/jViWY8SfkyxouFCE0avIjeF8WGdT0LvMIrI0NQAHfyW0Ptmvz0w9OWWDt1pSQEdzITprHDaSeL
t9St403XMeFnyxDZH/sjavAe+ZgTBJx55pWgW0xtcCL9a0BLDwmWuXur/u+EzpfzkzrkZUUwSbEu
RqLYOhtDsvJjUAlMq7NLmJPpMCq8iSABjyuMTJyZZvvTaD2jJEdgEg/QWp6vgk3ybcKGdr/wWTro
EVeaKPI8zzHfPw8Vx6nKeaYOeuqwB/7/UsM25g7veV6kDx2ePv89xG2KIADYWSmvuJsVkHz1jK8T
wogVkFHh9eaQVrHl8mKoECEV9JavEIofBxSswrV0NIsTw1xdO1NAhbDq+gq7i49FNsxsleCyi5Vh
cPt9l50zfighyGxSLBF/xkQz+LK6S/EG7b0FX1ltX0waXqMKNBuOvQccvnAvjXYdQv7ACPh2QDwp
8aOi1Gink2S07Ok2CInbwrGr5zOCobpw9JB+0zNg1OXT6YxiJ4CppeVUrcNsdQzMDROfdFA/QZdI
OihR0bdugF3Iy8sKfQHZqrK45qWMYt+CvHuOUnjCGb7D0PvahaIx3tAzd7/ametIunuAfW9sGH7Y
GUjUuqT3yh9GRqJ8LlOuWY0JCXyxCc6zpoOBRJ74bCAxS6SF24cRBPZqMQk3XFKO4hL95xGmcaF+
W2mByMe6VUnDs8xy4WOa/kx/N7bsHPSW+PnvL5SQO+QFBKDZ7ciJgRoUJyokDutMiBVj+mP+/7we
uaLHQkN3DR4qUsqwB8bq7v+i4r0LjcjuE2XahOb0tCE+rnrZ9zx4PNy23ZkFejpKc5w1drKUYfe9
DFzk2kXPRsnAWimaZS9ZyHBuq/4yog9CeUTBWdewB7J7qNcfDQaVbeLggob15r73AJVwDIWdZofQ
MNbQQ6TY6M2PXV/aB6/49W2f0d76P96W562SmGdS32ggXWUp2Mj6GMIIo9gcxQG6nVNdf4kZLYIh
wUtkZWb8D0z6bdqQLELy5+KGvjYkB6gVvHW3jthUOOD1RIU1K2QanSige+DZ1hdZqoa2mFE5i52W
52+AhRVRcHRPSHGSdKRCqLiY9raqb9QO9EHktbrmThU0PUniyrMIaPTm9+K1kip4kYg5k5V+HqlO
TuAop68Tskwu3RnCHl6N4rCBPCPRnOlg14PyjVVsY5W06AtHOaP7w7g0X4cxCRpT7VpNhsIniyKS
nLVXf6siI1LEg4pgFIPIxQy9StQIp11VgaMZrR1XHmBFfxsixVZTo6uVMoF3LmfB05q7t84kUY2F
Q/Z1E4UKTzX022mVsfHBUGAszxS/FjVtxMkQhwZmnxwcvzn3nXjwqjQjcLpjcwcUk6FZZuZBAEb7
Y9ASg4yPGBXX+sXB/qwIfNIMJVXKQSgY1V4JPV5BZHXeg1L6SB3XOxVM96LF+UkCYZ40dkh/nk7R
S97mH1EJYPX9flqjR/f1f9gWXJS398KXCW9IvYx7xQAaEzLIb0qicIVxGjffca0F4KNGgPJtmsdU
LJXsRJ1uj0lIN/xF8of4xV1kdBwSfrgJW4n6U/RqhbzPHduST76alMt8JR4LGuRDnwWtTux9e/uY
BJOQdK7Sb/zInVtPKGImkL8mzRnXADwFAj1tkyACULzz9VcdnZ8iLv4mduRZQscpIDO+tjAQRWiH
5RjhHRp4PGg3+guyiTX1oD2m57HUXICWns9JgbrBgzvDa90p0CrmaUlaoGR0m7y6CbHCFwjNGeQa
umiDsZDCfFO7iPNsecsl43h6hju1FOkvy6BqubdqrgLh/gEoREAlEhpAE7JfI/4ZJWJV95RAls/s
WopE5pEXvH+buy3R0gloyXZpbwHt/EKdLYzaN4ekZW5RIKlGH0E7hdQ1btXzFM4QQjNDKvTOY2fa
ECmeMjHyWruL/p52tAIcDgk7H9eJhcTRiXzuJsiB3Py1aUOmo37f/BpMsvGPXpWBzm89xMnKV4dc
YdA5mDCKjSusfHGlh4ds/WRx9WYtwJrZX44/O6W024d4Y6lAAuoLQ4RYXhwDYYbXQ6odMKWsWzfX
Tfx0q5z47EpfNAnOQRzSzBeAqX1lEU9DNBHDH7T18Ca1HHFwOMQqci632CCj3gPzT9Br+YH09OU/
4gg/7WxXGkUQrp080YxyzOoJGKgnBHcUWqVGe7mg6o1iloF8I53bRtIZH9OB3egJ9iwwsRsruuk5
SHwH5OoPMvBjJpzvSq9YSuqwVvsEytcXV/TKk56zW5zhHz3nj4ej7s8c35WAP+rf7qKzSmyzK8rT
wx5BGpvpTnPsnnQjxbrykFVrs6eNO2C4JyX8oAnHTZK2yETfXZItkOTDiJzxlIxeTMxMzd/1remb
VSBNyvoIfo+UbDcdxDr1AGUuFeoSsz7oiiLy6a9OcJ/0imw4ZE3P1D1V1ODTqJO6oZlC6F6wtllD
2Dl41lV/0Ejtf+PHyAzcumG8lSizraFbyo+J0YSllg0vo6JMdAjbH1HptA/EqWtj1Lh+9o4ZGqfe
ZmzKPpCtYCBZtTfi4vO0L4U3Eud2DIO+zIZn+xqN4Qtbxy1kUd0VHStdYyZ7dnWr8pKoHdl2/hRm
kwf7xPW3x0JAtHAidjPpgkyhWOUzV7Csy3IXm1YzmDUUEuMd3iJhYvW0KwFJO8zUx5vVE4JbXQfj
cdsrl/tIZY4X73I30XkWa6zcSZyccRw+ds+S32kntyiss+BRV4MX4r8YsTfYyJ13m+kSoWGarnOJ
FlaJ4UsWAc3oeL+zw0F+C4vLWow4FDKm4BDbPMkUkuSxgmDTzfOUsH4PEJIm8U+SAO2HY/tTLNCy
LJrT10/IPSJYwTUSu0VJQKTiffwXlcRLso+cfxId3n9KzP6JyvXWfq36Qcx5BZfAtxBdj0jiAuuj
btctTv4MDf9IbtUXtLOVRmwVQZw8wse3bSvTo92rgxKgMhLfGsa6joXwVb8tjv03Zs24I1i7zb0D
ScCOYjvi8JalwmThjyFotP4M+MZnXu62nYvrXaaTdw745nMA2I5Wp1f+GBRVG41XsQEJzcGtuvKU
/a0xufFac3qUwUT/hVD5tidD7tnBN4AnKWIqCaVsuGaojylyP21smwNaLNvkYv3J7Wt0aKMOWPuj
quRfikFdQna3PKu8uZvpscn5K0Sahr3Boe1fbzoMAnYf48mrWfbj/PIKmBDr0fMujVhnyhawhWAf
oRHgSBpz0qgEDMJPjG8onwf2AVfVqLP7sMRs7mFMGlEiTO3hPvdqcYl62SQOOFXkF564+kMc+IFH
popwt3jJvtFDYne2wMlOvFdt6N9bx6liTyvd2+mH/5MA6bRXCK4q8tw5YzbosMbcw4QkyqoCJfC0
NkPWmPyGQI+QvS0A2PbwPqlxahuA8rcc5R6i9wJCJs/ctBQ3ZhHoQQMn4m7Uxwp/kCJbY2Vua0c8
z6n8pK9/IrtywBUnVDAac23lJYyI/TSnWog1mQ/zqDj0jwbFjXCc9WiOZuh1gMGR6pHmaDVEZgs0
VjR8gk3dw2doYMMUNZ+3ZA2SnR1ZG/8QMdzZ+2laZWKipmmqHws3K89KG0k9lHEJOVvaNLnLw9A0
LJMv/gFhxdBRGApiq/66ZPTouEYpYHQSD1iQokgRcwvS4fdnnZNVm5gepjKop45U62N07u/6PLK4
pZQtiwhymVhYd3ZDqkOjtC+jIeO04HTgxfaZTP9SsTcDspiElCEJbRhVnURqYzV2eo7cdZBg3Q/1
33rD3psWqOzUHUOpKxGtB8jhr61pDjcrJsvwdiCfnd9E9m/wByMImcK6hDd6BmT84IHl9aYQe6mX
rHCbkvBc8IwP0iVTOEdipNlUv9AenFVCqUmf/utF0E2WGCNjjvI7qm5JN+hqkQ6DQAWsSguKRB/Z
pgIcT359uWhG8oVVGeGRyOHZTzZjyrarzVVAGSlu/i7Ij/JR7UxLOFjjD+KPvdq40PcY1zaDeRLf
JpnxpryPkCCAm13XbDOIIJ1+Z6oBl94bixd3raOjnsUu8ZhfZfZLp2Z5hI0oRzUDiatTxZpX5XAF
goUIsDYiRGej/rj8yXdpjKkquYBNGxOGEC9gPuU1OPhxXCpJY3RcSXKVF13oZ4dDVB/40WUUce8j
0CXMofZorgN4rp7zxSPXuIp16lf87HX0SsmvM26k+IKGbdpzugvvWROs0r0YNmSTVllpgUrUlcxT
GTrEVvOzxA2Whj0/m2PDyJvKd1aEB9HD7XHDeNZxNDdahc+8QnchuPAd0xfACI6OLC0z2svKVGmK
Ua/7DeTLM2mLgp69PHbwjb5RFRlPp79rmtVjGPM/j0QY9LkGpcykELknO7Fub+oHtsxMOEFwFBBN
Z/9Pjw2dojNJ8Itf2MvZB0+MiAYlukluSS6BxLSGk5TCSSFF2NsPF6BRVHaFIxoTLWy4/lDDrRS8
lNuSyiJFSeZEvus//ZvAXm38eEbnbmpAD0XCTbjMIodKUi5cCBOkj4MZPKSLCdFgwj6RF6w4ZgQR
SB+G9XtO4pghkoA1w+9dKEdvbfoHkbIaOCJYou6Et9ZYsuuaXA+L9mpzP0nXmmRO249BzMjNdKhe
dJcQndiM7eihgJHwLRRcs3bQeP7tq1hKaunoR2sNZaNpC/VnEi0Fic91eYRRhsXMs28QXXWmnNrt
dRKSpLuba+SVsiZd0J7zzp5addOVoL9F2tKz/0Hjtc1U5xJuisYbUyJDA+xrTubPJ7+XWQv7FHp3
I5opiOaiEbaaIGkWvYzgkJtVHMrxiSH6oz62/BesN+nqHzCabI1868Ugil9wnxk6F/tylLB58FbF
gyXPZ0iY3e5ySp+9RFvGtQw5ICkdYoqyJUAGv5a3q8tWCtr/SOcQ+jr7KfddiobvUxSKuH/Krzj8
nBuX4q2LRAHsNtW6+5HkOiEU0O5nksbFjoFjMPeJifLrqazXj8Tg7W/NHlsSfGTKbLA9g5/pva2H
flcxrqqINxnWONX4wS3gAWrdZ851vcYGopAwuo0NOTNxAnA+g6aFWcyRrNunFfMDTDRgVdapMlFW
r81pomyhVjK5N/zMxrFD2V7rk8VwcM/XPYEhqBjuAVOjhaEJ43ExFApPFYmcvv7bzAAew+GMzgfT
pXerKx1nsgXFZSZQ7xtUinW0Mv1nEVRaxVMKzSoY3Ez7KhQ1Za9kECN/J946TYANOmPjP+p6gJ0D
Zm53thto0X4u2fjPypZvSz9kqIo1pHjIqCBworF6R82x4qdla5zu2KwEN7HT7vJPrq1p9gZk0xa+
mZAXtJOAts3vpVbUYUMf2F4a4eIy8Fzf+wy+XVSnZ+Xdm3s1C0mKp0kaq98+If+eKpcS4Hnw9rY4
U3rIChEhGDdPjLldg9YYzxje5wPcy1mcGK3I9vmSvhLAT/hkFlXLb4aSy0o0qQ4xKqgx4dsH+jvt
QBlpU6ylJTYM433fE4NySjVHWecs54Utw6zaRv3SKsz2WSHci+1doow8mP7yE7EhEOBbVX7eTB+i
NK9wmvNAKwLbFBPEyBMXwAjrm9rAixijmKJ0OXWttPHa6wyhLOH3/QWYF5fTRXEJ0q61hUpz2DqC
cCAMHVrwPUVcHWq98n1usD2+v2FyXM3O+aUZJk+KiYXNEQKBnCs5eMA1aZmx07UvDm6bQ2oYi8+D
HraCdbNdG5D5NmTOQN62PUJTFujFcO0ikqbH17AWKs6+YxosDt+YsbJjl8ikBFMzVjL16QqEpUm4
2wCq80xgWBCal2UJI9M8ht1Hk6zudOUwk32SjZmVDUs73gmTdvNt4MeDrz3Mamys5LrAGDMMSFCk
VuLlh5BQydpHemJvzLmtW6tFrZ0aXpQ3XNOzznAV9EuxEPG0OMps0chdWDbgl5yIlrZ2BDYYzV2/
DAI1IoUNb+/VdAD3mjzBln/xHDV99gbgnXXLM+lUI6h3lsvkOLw3PecO9hq+vM6VrAD7jPgsZJnI
JTGT64K1nynZMM5mRIKS16f/vu8aQmZpjO9iUQ2y6xaLZ0EleIymmLRtc0+aloU5MeSVambsASb5
HJscloiNOfendw9Nuo1BHrq9K9kg2RknO5L3Ogmac92vDBCvVnCNhPFFTLr2nLv8ds5T+JSO89Xw
cYYkSd3dwbUdCI6+RfEUdNFfUQWuVjgh0Cipf8u80KFV1UPnOk9bDMhcRP7QLMS6juid0+EpRy2l
WH4FOW+WjXhWNkH/SzEUWVN4/O4BKZC1JbKd3bFNW2Ez7fdfC/YaebHleiw69rKXvplOTfpwzdtH
rjrYINAx5YfTNyKgZhZTqnwlglnrTq0Yy3T62Tu4anTM7Ez8eSlXj3r+/4b8XIF8aLxKae6wsFxB
UvsccgHKHtGddx211/XD+yuabs/T3j5QQ8q1J90tj4ptM5RvFXFd7WmFPO8n5QnvzSthj9f7y4kB
pfnyYut2ydcBJ/IuCpaNnwy1OxqruM+WIQ1NTd6xPgTM94Tp5cpIOm1/a1DnMXRgipt5sb/AAEy5
W1GMUe8+DJwDyC5f4EYwMSIYeJ15YaBVlQFK50QsuswbjdfihLqlITXavwkyR/Tj1l3RBADp2CFo
kch4ujGAzj2ubkJbKLRgdTTPbmz4IdkEnQ3MJwL9XZ1ntFAtyP9K8a0G35mOIpRnKKxuJLKCB8Tv
dmH+/GBFpXwlOM4q4q7TVc5fFAUYaRKiCHE+3yH4dU7JsT2/AXk7nIR7MN+KDTnnuXpXa89ieTI8
R65j3DGJt6Gp8ao4UH2sFWYn/dJ+4bCvD0SCAbu3KGOUx5R6lJoBT4q8k0UuRLEJV/ZLN8KOe1B3
8A6iN4k4Wg+/pHaYwqlaJuRYG1d0lkfEyKeFfXMnrvIS2aDonIEWGEeujAXUTM473f8xXkSj+Z8Q
NmUdCM4qo298NJu1AyJ1LMVVuexwuD10sTxTbk/2CQdhqfJ9lxYaGqbhFL5mvpY687t0a6RepCES
huqv3Wi+DAWS9BsYmrM5ZicgIYBBstf/miDHWhJODWoMO6l0IIPCFJoIvhbRmaeStPc4ES0c1lhT
oHeOKq5w8rPRVTA/Xct9O1dZx1k4a5WmUd6g8ZSAfYk8+GRIEeVdowFYo1R0y5xkH0ZTdHjzbDcU
mVE+3TJ0Rq/I85mpG6FzqjhGIklyiIveSxvXBpLD/rjxFqhVNbvGOZvJlBRYg1khPjVhncFPZLb4
SvF0DjZWlTgSd07Zz0w3awuje72MHaSfy7LiRlHFNb5m7nioiWT56W3jKkyo32Ni1o069E/B2iXD
ILzLkzI59A5S9bbUuEzitOWHhRwLVHB881t2O8UINZTtsx5LlEIXt3N+1oDIEzAWla3MBh+JDxay
acnSPY0wibpIuOLozEbmGRBoPco4nAhG/iBRFBnp3t8snln7chM1500Hx4KYmXFoCZh78m1GA3AU
X70ke7imL6WAnOv+IRnopZ3D4WQGP5OyMJUXy0PeiYoSr3dnLcGksD/LGhPicXqxrF4uBoNg0XfJ
Q5TAfyK0xLmaaGXVGyST6KsmNyptb0VdcBGhOx/PdeH16bLQMZl1EuVP0uNuZ15XR0r2fWhR1jAk
Pu4AXk1qjVoDjCTKb+Ty9r0QFfpssJszu1wj4/VmdD/UEJqcZxy0NxUHBt+InCihrxn6EI8Q/bUx
yEZdKgF0SHR7djn5ohTO3q499ufApBnEACcq0bTAefBSUzzLSXwKQPEVReR4hE8LkICeAHeEqkcx
d101ty7M1YG6ixllso2hcWWmYHdcUi7yLAkPUDtrUWf+76z9NmyWFgd5EXnn+14zfEIHarN0EjBm
/iv1whtDD7Lvt3qz5qs+FjTJCvqhz8cbtioiifjy3rqNsDA5abrl2DeDKj5DdnARpjDp81r1TzE1
v11s9Zy4aTELy9q4CUwEykYtJSmw1zYohuGJOHptShcXmEYDiK+UePNsibtviZ18cgywangSMBxD
5+qrgU42kM6vhHYnfVaiXgRnLs0SXzamqgBRLEeuTnEXspqCd5zIEHaDzU6by+cx9/293wJc3rfq
g03rgsxxSZi+YhJYWcn5HQIbhUb8DAsFwE5xAvQ0RWDfPxQEk1ShAz8vZZPGEugC9A/129ZEReF3
cN0Nv1NxlIZruxQBugMkiSJJaNe+jZ1eSCBfEOgRSgDvIaCpZW476RQbKFLX4+9PAhG7o8TIqBRU
GaEHSgI+aVKtG5lktGkcg9NrMoPnl/ksMOXqhxEllyy/fU3IJkZnbSn1e79jTBDNN876MX9IqLpj
IxTwPLL1YVOrYXyi5+adiuT/FGcSdporOBbAh8dyaCNJqhqUe1MU+C2d8HJD1wfv0Hws68mlynjU
JALtzLHl1MJPZjoNFA+GcCAAwdV1/jEB4m/85nlw58a3wMBjprQBST2JC+Iy5Eayv82KKSHsj/tK
QQItlHKQXj89B/x+fT+S7KNSFo1ebGOJpNt1pdjXea+LGPrsk9LwVCej1IHqhGfgwufnTrtrXln7
g4NgDjSXRpWTcHA1MGyOE2MEsn9pJILurxwvlVxlsvL7LgHxeBAG08PjRGEzqro4nO4pdczbuupx
cTs9E1g1wF4WhBl0hQgolMMBgvhlXHSMXfFqnI+cypI2mcuHzRoxyoTMJDmez1j8aODDse94Wrv8
TM7x0/ja1JICOPqvFwJ8S1i+3l81Q0Ps5X9uI33tOyWd5OhGGyvWJnEpXZbXjdcSRJNa3imtVhzI
bbHLOJNNHHzlJu60T9QWFPVO/5OcxdYgj6zFbhHPIFbWmaMDcPyy9PKI10yziTZjW/G65Wl1DYg/
ZQWUkN08FtlY1V6OT2V6bX26mHNwqrBUz2eqo9Echze/Ka65Q452X++8R2kE4lDQW/Kry+n5BA26
PzqcWX4zC+tGL9PUhaVNC0SdIAP6ub1hpDDl5QEY4J+oDYpXNaxvbimvd0qIWfBzvZNc8qOB0hgA
FMZAyUAPGPsFgQtLIpdT/psQJp6ZSBAcgkOZNPJdw+I2bZQGk/8YfdSgC5l9N9IBRMHWOzCFoPDi
AJ1SQOjHMYfkX3k2zH8nqzWjerXPQFI8swAWKvkEUHLBCV/ja5L0+2MLlTwOJsr7bgDEjD3c1Qv9
Uv+28+1z8oh9OqlbLO9ecmLpzKV+tEQGkPD9Qx9beb/jzRmgdJApnrnZxwrNijbGYOR94y1dNkr4
8UBugabNfiqulcv6UP/baxnMFFpd0xp+xNL87Gf5nKkjHeaYsawPlV9Xwp0iPPf9Ux2wpE0Ld3D1
ZyL3xSSke4GWLerSBCSl3iJD+Ib+Xc2lqjDbppHf1mls7D5SB/sOymVP3DHi4xCZ+bwi+bFumxSX
GLyT9gDA9y9BaopstogXHTESqDXocMio0vi30FUDitKvP/M4dUqeCxlRhZM9U5Smgp1eud38ZCm5
mvs7tXQYteVQk+m1+KyxEnTI6iuMlSbdzIgk6XD5NiEnCTetOEuKyEpyD7GDKHlWnI1/M46WX2CY
J8tsaqfLytMN0GKICPtYrUBxQlq+WieOho/W/QEv4j5F2VjijtLPMi3BkobCwSZMRs++TuSE6cy3
mG2LN3lBao16JlcO/XU43sccK/4s9qkduZTPksp23DD0NCBUIk+dXkhl7et5CKMRZkdCFdBuMFZO
4g2NFOfMAF2VDt80zHYsbS+zx/fogN3WC1uRzqEwM4xhDbN84oXz5Jv772FJ8KOgJBjT3oLlBkT2
tfkdx6fDhXFL+DHBz+2sbGeAykmvULuYifwL8f5fNVdWOpHC9Br4fHqo+lR3zJhS2zbyKEo8RKao
xtGIlsJ4Idze+hWEQo/JymtKbcYdDeXYcXRvu/tREN6rvMbHQlTI5tK8WaUsO6JVVL40sQrCv8b9
IeLP3sihBIsbjWDZ64yjlp7otQZeLHlkuMfY0LCDz0UOC2FkISm677LL0nV9vxKA6/VjlhZr1gMA
01xb8zN7BCRHCkP1c5g5/7+Rj7K4KXk++vjLdCln4fE+Cx5dxvLyUA/H1CnmXvyYjptKuH/3ixU6
zw/PnnhFEhQHw8oeYrWsPnsiyYmcYbr1KXfYVJ9yQ/ydnF9qnYLUdZ0AA9VAlUxm/lHKQsJvctOr
xRuZW0FUjhR4Xxj8ChoeaQ21ANX9IO4CsP08v+xgAJ0bf7i5l1JGpEt+9LTjXlgqkxXlWO9C3a0E
VFssonJBE+WJAYhmIRBTb1PVPyspkJiLp5jiyjvz/UQPNlBBUpmdR09gx5zKi3HtKlY/RW5IICqh
11GhZ227x/lDI5shBg27IiyXP3c5NBizQk96E+DlKCMsJ/nn9ATnG6Uy7HcLXlxVD5eZvCF6m9Db
rb2jhiK31oHzR1Dd68DYOCZxgL1XSRubW7ty32WKu6srhLujVzZQFZTWyllgiQ1PHELTPh5D8AAM
x+RmfCE8jIi3XA/qHJtr/krlk66xZXskwP2YMgv2eFAwYmBjuegbSBqUkUUxYT49FUlZc9ojQdgJ
wtAvo/80+K6yMF8+nsFnmpnauJjWeWyX4yZIgB5k2oxVqxcMFuRmQi69EveY5k6fswhuPHTiUSH4
q2nOVftn6AYiZOFaZkYAnSLd57Id3V6tGDiq2GNm1YdJSZ252cJi8C9NeVIDeDNpg7esOSbYDsOB
nR1iJNbZVFXCA7RHaVoPt44kRtwP+Vh+dLUnliw5IN1LkWASUl4X/K+Gz1/olh835dKS3vv5i2Lo
neBAM88j79ahBXXQiteLwsJ4dJ7Zs+mBGhntrgAHvY3M5rel6nNCD9hJ48VOY63bBEQrFZipFg07
5fdtvKrq5OgHdunv6ufUOm4G9QjBlWF/4KcqDZvWheS4+0JCwZLDaBO+1BSvuITWst5z/0pqVMf8
s0DXOsN8e5nyMfBh6DbVHnS9lKP6bt/kWHM0ygl+mLVyR7CGEDNrcFQhKb7SQHHIN7xS7KZLtrh4
HD12/RLIckGOWGrgKEZHmhpABAPXNRZvHjMr/g0bajvST1dLhxixw+fWwmzaCg0VkHXEKyg1pR+u
71Ik6GlCuhujbN1NOcIe0hVHtqhrzrUm2cigfSBZgIYmknHqKiPnm38+eDGEasQa0wZRgXVgB4Xt
i/AAlSprDCE8jvQsnGjwXk3jJXKKgNFso7Uhlm9joms12Wp1gNLeDyjdesTaLeFFQRwBNOBMzUr0
RHaYLyuGnSse3ntbjz6IO3yBkZIqGGdi46Iep+lTrKzNNxADYzSSoFwsj0PMjGLpm61P1t2q0/sG
YZMuAKwAOzlNfH3UVA8yraNYFuaeYvGRaX4BCVB1fSxl6n8ccJ+FY9qm5+rgEyXphpikYCIQGVLg
zzD1RlskMjl70lEcYBbVOHY2cHdtXjyiP83em+TouYLwXc7HvokOjjEXjdsrE5r4DESfFMqngnQi
alEEw+u3Qe3XNN9SqkA+eV4h+/aMzz1ULRNYSbTgTgUkU8w8Rt1XTozVrlB6OKTUR6iC/Z/i1gKX
DIPgETK4wzQuCMrLsYtWi+voVO/bogaRgnpqmyPvbEVKdYWAW3oPO5993r3YBvEhBCQ5K/h13MgL
WZJvIfWXJgyD6f52MrI7IK7L6wkwfijvtcb1Wly+Bi1JGaR+UfMKHfwNaUkVNiGO/TbyEH5O2yET
tALJNQdvW89EDJZJB9kTrtAhlMdFOyNg03GSACHK05/jxmGvn51/lr86GyEGbu1PAgKbuRvrkdjt
F0ClB7+tZfToQo8t+KZ9PzZIFUO8GrgqYgxHThHEDkgie0MI3En8WYE5Q6dlp5fCApSvrb79JA6V
0qe8Z0bOMWQgdRs4T1jlXZ/6sXri4r1FnvowC/ZJvkkV52QIbbKdyC/HeaqvrXLbOZxZ+CKUggBS
kE/x7ra2o7/W+d2vi8nwrp9LQ40RMhOKG+nr7ENvNMjxEP9omdR5ySk1n1BiIPMOYjq2U+6su+cJ
MYktC47pJIfujBMLLrqsJvxBbKrPPWcywBD+CDi8lOyTUL0ims3+P49Fs4cJ8DO1f1/oe1h37QS1
ct08RNpc6Zp3v1fBzuQ1Pwf54nJX+Cgbyav1t/r3dT5sfKD3cVvMOnKg/1z1gLB0nq/v6SDQu2+p
viAO/MHV8AdFop/YnBJZwvADr7NAR0j5J7srS8lELXOPkZq7PuhDDcE8gRsg63dhV4XmbPGEbATT
M3jnp05B5ScHq7ZxXst5u91MHCeiL3MMqH878qKuNCTeml9Eiyu8mGHUWFYJA+BVMnqWjCOEc0oY
M5CI6/Yk0avot7OlQSY+wmuTMhfUb8TyiFW2sBP4pr4wAF18EUSATZfKMNGfpvJLDlkMM9rgva8R
+D3fOJ1kAz0BGvXXRi5A4JupOUfoxoWSlqAaCPAf463qjRSvPJD08661/VOB3KlhzcPPvHwf3GTo
Avs3TQwux8EJgpacuvAKfBuuqF31VCiPUVW4rkG6l91pPa6fWt9UdOnxuFtDZxWprQ4Jeary2+5v
mhyB/rt814FrOeeyAMoDHojnaK9fo6lzv9TEa97H7WQxer8lpMIyEHJ+0VbGVtFSoqmszrTYa5zl
FDP+smu21DkF2+eojNEqvDb4Uuu2xqIrwjmGI7Oi6Ky34NqLU87l4Ws9/3SnncquPMaY0wW7pXsJ
uuJFRIJ2ReqH3DcBkwJHjgcjxSjtJ1aF1m4exxW/SWDs79kFPAFWdlcHUbUNkzr+igTrum6fXPCZ
FOWJx83cQaW0m/M1kIkTBRzzeu+2mtqF1frJP2czoAcpe1lUpzsDJaDzpqrgx3of7h8/GyjjwXAJ
XtiygCP0YX2Ny/O9WxgFhDTGGQGnee6HPIThQRYoQ+HKO542nOIeKSGCHA3eWhxK31roQXlTCqFZ
PSdzOjakCo13qWAJD6HKwA2ClgJxV+ytXeciT/P5VmRSCKupnZo6ZjWlj0DXT+XFM0GMLo8pmN5y
205iNcoA5pxq3dtrBtY8r58L1+Fj+9tnbB2LqxVO0GbS8aKnT+2LNIan3Mu3E4dTOLJLQjXsWvaI
I0JrpvbyQyEdDYOX/6TEpu/JHdEzGgfkDrnpmsaNBX0qeMn3Do+YyejzvrFz8M8BmCo02kvDWn5c
r2MnbmokBsiMYUWl6KYLLQJYonLWOi9I8UZvOurFtcg9T9CY61+uiDVh4iHDLrbTh2yg+Gtw/8Aq
HGa/8G+rrDP0pypE7jM91j2H64CFZaLbrJLxNdsh/Fdl+nMTo3VvnrZ/Qc7Zpvgx87fEwi/BENpM
7MR4pYxq1bUyQ7hnjqAxd4szqjF6KhFtFxN4IUjJKZ5h+RDL7+2/Mr1higLifJuC1tJECrJQ2/vn
rJbYhG+4Sp058y7nJx887XgWHJkRIscD9SPKhNOdtEXBmZOd+AtruOju+RkkIZwR0CxzyNFhRyj9
btuHNlDZNNOQrmVOrt2qnqRrQqbq2xOk8UxRnpGJXkqDhquJgpVArDvif9DRd/g6oYUchVoglPvR
kI3qjHycpcIMNWsz+tHvQxFc9NB6ZrwGIKo/qWUt40yTVDpg3hCfMTuXx0as7f0MuuEGNMYW01Df
h2RlIP0XzZSNgqpyNh0RyP0mBKDGurm0ZuDpPcdSLhOh0Oz0eDYScTlITNbBkB9ZKHyxNQEKG1Sz
vuOmv+wE8aa6zNfqINRQhGsdgMXcyvROQeMFI3aLFAHWbFfrNmuSpS9I1bLcH59skMck9rjnQl+g
80tuI/pkTxwRcxu+mwqsvy1XbyQuJCK11ZlbzIeNbAnVTuOKNWAGnknAfwFn+IBMRoQvKoMWLVES
ITAKh8Yw7ZwWN6tI+gPTGlDCZmBI92UZbbBiv9p0SZI60ojw2uOor8OE0CpBPqkvYpvRiolXZsrg
IFU2m2gEPVZHbUC6zI7D9Yu9jWgk9y4sJKvlSUmLdLdob1ZSp6piqKUF1mjFe0Rs3juEX7Fhv01Q
5P26TTTZGuo1tDofCMCQzSszwHPht9I0M1k5Qw/XqU53Llc7vz/6lcRvlGIOdPOTj02paQc6Na3X
9Kn8U/0bOWWPcXhX0cvoFMenqbTIT8TAjW3A7OuvBNX2OLxPXA28Qs8h+5GNri2S75GQpm6hH/DF
sjMFLKXx5y+1GblEjEU3u9iBn2dSWlcigxE0uSSQlBZBV9LpO2bB2XYBkGftLAIpgqderxCxEb2d
gD3MFC9kPU0rZ09Lu1ZJOUkRsJ60Hni7v2Tw4lMEhBQJo3KEg/Z0WrXkqkYrbI7NwgAs12kA9pz0
SnNxFGZm9xEcunhEKhzfg2jVKFCTm0Qa1jXE8fLqKR3qGp5E4InRIsGQJUA8j5ihWLCNlUatBvrF
xvqqaEsd9LY33ZJVtJnxTabDmy7q3NOifuRvxtrLl/Konjz/0w1ghRT0lLUDveMmFleGsDdFwPh6
eKEQHEx3xxf2hD93/g4xVX9puz6+2/+ZVbWrl49Tdtaegr0clYrMeNz2t1/zVDibgYpw5KYwgR5w
YO81cQig3RY+EUhF+y46suNkzjREZbttl8GcMaKJM/lLEvi9p0CSjSqaxrOwyqCIWmAM2FS2R+Wf
Pj2KFV3I4kLlm8ZfdBlAgbdu3rq/86x8IGLVyHPGs4V8F/C1mS+6p6K55yiRfQVKD0v0MiVR5X6w
1HzF8uAjOiOjT5oBygtbZ6EWZwo4UtmYMQautltMWjL2gE5y825X/kyupb26ycIN3u2778rIDLLa
Ivg+bqw2iGcFWNR2kSBw4fVW9vbHqEUeQRMTcI3IcQGL32hh6PKbJiYw3a5xU8HGyby5ULKkljj/
HQK0oXD41kp3OHJLeObx1K1qDEIkUfnZ/Lou8ga5oFrypT9P9ixTxGbeVvDPzjlbi0RPeZK4gwiY
CbwZcW4l3i3az6gLUzLAr2bFWoUCjaV7yIypHTplpXvzfu9GY2sA6bxqm1YKr55emPl+hkx3RG0Q
xOwJNeluz+DuQnZe7QHmRJFQ9YV+tgg37rOapOWW0FnQeCxQuFNfSYb5n2HPXhHbNkhjT2LKKn55
LMSBcvUDz69qaci1cYnAAN0T5mxmgs4RlCguqY0X/qlKle4Q6uNrEDtBtRPxv/GLHr66MDuZaK5I
WHIEq0gy/WqO+Xwy70EDOyKGkbDxJU7BnWdTWjWSbo+zTiVG5Uhgb1i04x8GKE+6hGFlfhJPeANl
LpEhjgoOwJo2TzSIP1rOYVyHmMorUE+UCL/gylzv99dx1a3dTSOsqtDAnAMQ3OVPKtnWd39WbQh4
Qw40GBRHhJysOLZx2uVRjGpb6bdj+dP0zginlSP47j1zNjehb7+wt+ygZLT4Lkar1P142Gx3l9oL
VWA55SjmLO0S5iicZWl3CA5EjbSZQsYSDAlLfsa9VuFuGytqKYrJ+DIdY0q4nQFbJ8ddOTsCN2mv
4FPsv5B56PzyGZ99KuvoF+hY6Q61jI0+TQ5NYDez/CNPJp97fSGrzijHC+nDeh4Xn84KHtRNL0Q7
7QSR2uHUJ+2cGAuzHFvwG7CjRax69KQab5w2b0YdvnF/is40CfIrnLJMK4+C/Od0MyjDPwd8aWMQ
EK/0qdBzJQcn2P5gpPy+ee1/OdYwv6uUZKMEYSWEgeV0CDLR5a/906hnVWZWvC+vXr2Ca3AeEm/H
GD7JgrSXynesn2YCx2CzYWYROz+FaXwQEhD6q2GBG7WclECLK2eRomqTgKPVia2tKkTeZsjMi3lP
1i4kDsEYCsWs2vTx9XaullS1fLyJSlvgg/G7BsifgkEH3xEqaKiBbubHnwet5j5+pks75FTyaLL0
EjbUvHmjNdi9XsPPtKTNVzNo7vreoKHltnPBQ3UWq+Q3kaVpHhiJzETTa8CQ1RpH8XycFNj/ZebH
UlA6P0d+mHngm9yqjYbQYvJh7DI8B4QQAfrQdebPbh2+w5z7lbe13SVTF23wmI8OKpbvude2b0iY
m/0Q4fLXMrq2OY6DB5sgBgtv9lhvpSCt8TGyQew6QWwR1/VNzQZaSROA0CSuyZNQLOSR9wWVdDnu
p1xVQ65GvI3XTzydHwXI/nHBPvDO7cxNEZ8FCwi7bxeiDXyw3fze5d2q3nXiNP5xvJIyMO6BH9fi
Y9+vrPpRm4BIucLQG5Nx/GTfPFkhOC1fAg/GTApcaJk/Fj/hCgqe4jwD/g75D5f8MF8ri9uKSnA2
UrG1sjikglJPW22wBzDO7gIlivELqmfy4of+8fhxh/Fvl7xr/8xC+jkoMZ1IN2HYTOjpXsvVQF3O
LsfT9CFVL/hDZLmjIHEDpl4m8f9yOtI8W9+1O9s71rkIqOQhuLWAuJ4v2RJKXBg27RThjvKrf7Yw
4NrqzjL9TOPm0TyubBJX2qlanYTX06Kqeu2OH/nqxZiVNJDDepPb4912PokyWUiCa+gO7bqILLBA
oWqvrikpKW/+9CIlOVmmNA+6ik8+7f+RjnUD1ilz/mTUOFRlUxpyeerZGWHendgNFsvoEssnHi+7
W0d6kgZ1VL4SSNnJZDNELl/c/cy+1/ofyUtHcJSPEFpdgTZ2iK7BE6j6g0OnNsUIAoOfpLih0rSy
0u4taTHzxOxrsHWtKMz2ahOtBbxg8TKxDG9QAt7SJMn+9GFLKLUTg98pfIbhb5kbbTasqQgaZ7SC
A0D+sgjDLfeoI7FGLhpOplIkbC37jcUbvfivAeofEuv50Oy4GtPQfza9ytQyvQDCawt3l6Nm107F
SJmaZ56HOeLjsv7VOwwcUugbTRKtsaUUuHoRzY1ER/WXqx0CiK8M8wdO9aMPuuIiiTlZ/+086kz6
h+daFiJv4bjyqyQ2Dh6iorW5bcz47H5MueHbHcv2E/WfLIRwEH2XqOqBcm3Gyhr8xwfrcDt9A78+
mo3vmrboiXv5BtDNahHGQIzM5SRJP7x1owIBx+amuul1bhiwBrw/5T/UgbJ1WEQSNHTN9X+UO+zq
S0Avv+Ff+CgVe4O3M0omo5v8GQFD9zvPgj86fYrL19vOiw4ePFduXlYpKmTGvVByIvB5+6LjBkDp
2dXy0vDFL2/Mr6E5V+DHQcXBqHRX8mRoungumhgPGUoKz8xbNQTF8amF8hJXk814ZGNolSld7Z9y
0tT1JN+3Xsc5ipvxT1LLoey0Y+CW+TqryKyEbSoSUn9gX66w6iKXzymRy6YwfzK4PeOzGgfiJib6
7ElK3I11s5POEfE+QRCk5NhqiqmJkfYna/Zh4eYDUiWjYbP4LL7o8RxsV+0YfUVGrLaDrFx9+Pvw
pxOrFbGtVTcaupY7+nBOsvYq1TnrsCUk7gPececalSlblyAF81FjTvo936SrWVC8C4Nn2S/BeiXk
YVERvrdpbxUub5XH32fJ6c4r2LGSmsfTAT3jN10LsO/c/vI0JkdzQM/19J3RQZRoPuaI8LY863dI
xCPmCz6sJ6zQqWqH8WgWdUQc3y48LaBhYYj0eRpeMDCYwuqhbsTL05RYDvhShqVR+BYp5d2J70l2
4ssSkomIrmoWjxK48iZMzkl3x3n7pvIIqH+7lMhJyijH3lNDVMZUONGXRN0HiME5qctRck5F3npg
rdEByEnjdllc+ZWDmeTOQ06xVdTAy7TK8HzaH4yCbiHLo6bmDv1xHZmRb1S/7J9LkQ64qOABYgCQ
/sPia83/vSbuLmpAcGYqZG1TfuQFG5KCAddJubOutwMfX9au98UEMtIlVQ5HqFw9c7GzJDKp/TSo
LMHVeSM0BFN+ZH2BA5vnA1Cixd9k/NEmBnnZIf1/VTfla3jWFlifm+0UyGq7zHDi5oDbziQowiVj
J4/Dl1FZk/rPK90hf8UXbrsLHqCExmhlV207n4DsIw6nQPVZEsFdiikYirv1JglTJAx80vnWuma0
oQQqh5mVkvzy2i4qE75yIfTXfTFOJRxsTY/bUDDTc0KGqOOe1h6YQUgmH0l6tl1g6mwouf1zZGip
xNdax6w0P44MPSvHHdXkw0hFIYRXOmE5oZ1HpYNTv0K8E7MBohdTIssaDdVV5RKSFWzAmfNTlOl0
32ozDtonDHrMdzIv3cvvBsCbVByazdgGL6jZFY2BYXAgynHvZKHy2T3InGrnIlcLTreAgWvbTK/v
Eksw056IWNtU1QXftY9SanZ8zW3o8WBWTm1hd8CHaRGP0mK6gkfRU4L1ihs8JCTkJBpjMFb3B2WD
Bg3ufTwOBnZO0HFrX4F8ipiScQh6vMiVcBFGEHE4yZwjca6tJjFVltlLpCKgjSHZqiSVKGOQEW79
2NxJ6B9WMYrsCkDWg0XJMoI3N99IJCrHVPc/X1uKpBfGsjGccpAXrjs3DIt4HsMV+Q7DMGR+QcQA
I/8yQN5mu7LfzHfm65qA/DyfBDDIcH8Py5yReoZAx8wMJ8zy76Raq0BRsNfnyaktonmAjuWHwZhV
u31/IuapmAHI2lgPcFTqnKiQ5eyGMsmWC4Rkl0/NaKZ3is44iPYHZftBH+q1jaSVr4G0OJAiwrVw
T4/AKKDCz0HVYPhlIiF3RrVw6odlg+9uXrwI++gh1aSOQrZEETE2A7k10ZnDKWf1Deq6UMGz5HCl
G3hXanVmWIB1E/KV5cV1jfV63NiRMwvLnR0YdkbOEgcVmg35eWcWlv2aTcEHdLKsbNugxhpsvWS7
WCSxKBmqRY7J5dq4GdrCvGEeJmVSK9iCp7ILwwEvzc/D8aO4CKnT/zIoEZH78HQ8an2vwyA5JMPL
nTcuB+gGu302z2l2zL8HbExYZF3EbWjl+fw6RZvUPbpAugXrRE3QGN/MyglvYQK7JQrJhEZsePzC
2NE0IhBWmlDCgfEQFCl0RdqImSM59ebpLoJnNPn75fHeS8sJt/TxD4Fd5enm7qaP3EZw4jkfuz3z
hWXSalDwuN9iDYHRRbbEzqrKSEfCwPLAm+UlMX5ZZVSuzAEZYroBLwrkmYFIRtqd+im+P/gmAvju
z6NgxSwS748P7or8NIZdyRuv+aFAuoNfMVb57z05pXvY0MLqmFE5w0g9Fqu4Kz1U3LqzmRkMtXwY
jdC2mtymhwmiHzyHnTZrFtXN4RlDjZNDoRlFb9vv979BF2oONNNoikXgaGF4ArdrJPd8KHGzCH0B
PIHr6VJdWnQqV57sCHtwBADtLw5TLK2LfOoz6ak+/bf5E2ICbpRy/Jq1LCGYyVqA2ZT0ppqvfjMv
DTqTFaZcChLSZ5wKzR0nw/7/MzktU3M2ZdShLgaerbnzMqB2lWbpH+3GdesxWkyBmiGamzOcue3J
2EOmdooOf4MeR8ULIM4BdUOre7TPFoLyWd9LrlwpCEq+z6HsrAURbHUAe2AWyikjy8nYU1qFADQO
O/a5QDXAHt/Yr0i7yPuZA3XoM05uxFLexU31dtuXOstVLI9QLupEGdlgIb2ConRe6ZtSpMZdY9sB
FraPaB/OhaYZsY7j1KF2bCy60yyKow+J5kEKoG1tqZukuLYZrOkLEI0cuIY34cRc5un/Qx9ZN270
X8gufEfFP05KoZyH8hp+S8kPNuF4yLHA+ajiMd9YATy4hHaWCcysB7UH1X/3GaFsekJBii2qHBmv
PXsteQ+ffKtVW9yUpHRcvg+ht1THUYuVzLR4PLoeJjYhB+kK4KSAO+tYM7KOog5nZLOTSBjXpEIy
43sQCK1i+C6AWPU4/QhsMdAAEClZe5QfnUp3U2HK5TAv8K9yiOk9ZvJNvJF/98iFn5SAIjEh02jT
wWiW008bBAPkyysKfKAmlaDSSiEaTrFy6oZ9jesf1MKfAyTAAh+vZFJdDVJaQiBetkj2mBLaIYMf
VJxJ/IzOpTnQv9FbT6EBTWUjxU0uuKWuw4IusgyryjwPxNlE3/vznd3hh5cQX8FDEMyXZYBCPRiv
ASDebEQT0ep7FNWBzH+HkA0dUXNu4ZpuNFW4ezrJZCB9phVqQvVhj4DIguwFbI9yZcbcj+Nfbmwo
4HsE8xeAAhGXHVBShD/gvB9+Sw3xiIFyLGpcjaGfiGWI8lf1VMgTi6r3aPOSr2uGiIckPn3irq4R
O71z037P7i6zWhr7XMzFyJTm0JdZsYC0PfuFbt8wPx73bkxxGV0IGH7gZG56WaDOpzak/b0ABrnR
FnZGfE70jKktI10xA4uXo0V30aaiE/Qbe9bcod0wN4VPoW8oCQoIsprA0jRvJyrJ6md9FzcBgd46
Ed9lCuw/P+1bQnwmAxmKQaygWxsSY7mHuSEKM/+RmQ46+rRfd7ieWPz7H1coh4IFeuv+7vl/iGzV
XZAuS1xSOkH6+bQFemKkwt4pYtWjJ/6Rwx5JyUd5t0ipWr1YIqUCQxlFGoQXJsp7sK5wDHkxzkbo
+1+eN07Q8tqHGSTPid0Nw5g130bE3/weAz8hbxsZaHUS/J4RyNB/7dzE2NLaolRAuqN1XWfPANhc
Olq5SCHJdnuoS7oJovSR8NFUi/24Uue8LNnG0sFkXO0nRxOe9/DFgDxfuDXxthrwegmS0KpMG30N
WcKTkahQkUCKEZ4nkrgatYuPhiKoPISlSaDNMipTGD7jq5uRX4bm3nsUsjd5EOZly6Qy66vhb6GX
xIWv/EtCe5yqAe6NczDq7L0rCRP2XceM1PlFH+4gA9unnEbgVwCT+AMmzvjn+YzeOCPzcUD46saA
qXs57cxO0Ze6ZpMmJgfgfP9dwoQLs6bHlrh74Yzjs2kUYdNpsgJyYc4Z1kWFWWvuIiTHfYaH1wFT
Mh3FCUD0eZhIqGziO/UBUCHqJRHqrZ3sBbM+Qap167AyY6fzZrGshZ3WgQvnCwc1zMnmO8yt205k
ukwRKdllmFZvdra5x12DY0VH5K2buSnLw5TKL18a7Yyf+eMM7HK23tBkIe8hXFh5hBDN8o0s30Ix
b9gpwfMk73f2LsVW9URSmTTWkZ4L/fRdha2ZzGulwv5ZFG/JwZfMNXqHJPvDEIvOBYnMF85WZuUd
VZjF77fhNq3BfryuWVvSGqJiDN65mcpLGj57GDdC4EBCLoZ8ZndxjG1GLRHJHMcjQSOHf+Iho0/C
ifuK3NwhTwFwMIe61yEOYMT2xjkHxeaysW7HbIoW22lOo2/jnuUj75Ci94pVYsn1GCHx4dMGyad/
qbJo2XXyM0KJRL8+1aH5H5aNaZdoVAq9gDsZ1UPVam9zc3hl9aOV0ESrQV1agagP1I1MJpiugW6B
k8h+9wr8NUHMxOx73ov6dmrc/ds563eizOxUczqwq6IdIqeA3Q886HB62bA88qn+dhBXiwc2d6Mi
rAQ3gVJhpmgvxSj2gMl/wFktD2Hvt70/haeH/ZBMWCjM2AxMbye8MWDW5h8CYqSUD+opluct46lJ
5fBV4K+7VjbzndZYuM+m1Se+N1BieV4ywpdrBEM9B1V+uhyfqPL6GNzn+yPMF1o+O9Ef0fM1qhxj
+LG/cbPgdUAAmMbstkaXoNtThd17PdaB7HSmYwEhoB/tM1r5KyHWRt5R1SfWMzaMTnEg+jWP2+5A
rSY7q1uBZx/UKH3cRiyuEf+42Bt56ceVnoqhZztBZ9mearAQ5bjdhq0+VNIEhm45pwz2ht2jsa0P
c/OZsJNQTGN/6ZZgB/aAQPB+fioNxTAAnhDEyMM0L2tPpxcgYkWnAUHnrKupaIrHXFDvnS+cVLvq
ZEDWEba7Vzuvi3JkVJxdVCyonbQbEk65jWnsRx5/502bEfdvH/fEIzPhjJxOidoPv57XJlIyD/pi
KfW4lfRkc7hgp/PnMe0wEmNXuUL/1MBMWxz2jM9nrC1KxnNcqPrQs8dP5npMfihwcD48nlkDPnp+
HkCvEE+UCfyPdtMHRQmxnZIU4uAnb7SxDyVzflWZ9O0HwNF3TDHnlekIgTfckNQKPiM2fVv2xzce
byAJ/qQgEhTHfJrUKGMuswVQxT2d11x5DfaCht6qiTbE6NhKpJN10RSQR30XCkEergEKLktdRnh9
tG5QskwMiHPV89guwstQFO7Vgqre1DzbLzp7ZRCY73QTttL2W4Q30/xCAFknIQtiGGi1K0nvCOkb
QpIErs2YAeMp0ypwcml77P4c+5dqD+BqUqpdpH0q8JEryC3aG/Ghpo8udFjiydHpuBz6AV+xmu2k
p2weRWa1kNVB74S+H50jcm/r7uiljSEeEliq71cvOvWUQ/cP+PfwmHNe5Ecu96A9MalRf8Ni2JQx
dUZDGVLEW1TLUEz8rJnDLIq0QENvyXKvk2HZXGGcPVaQTaRPjVV0uvkvkCcBgF2bI7KE0+szKk1L
nTYsYYTjLIDId54m1jyLFca1eKvjRJ6UD8mzLBjjqicbo4KOMIWmDPKgJ7xmNlznPojrDRSgGnai
1tF9A3yYQMYOpa3cjPoAwlxMpk932XkNr10wgx4SumtTB9qdhQrsLC3uKiCxjaYohrJa9N4KMVek
7TicvqYCafGKz7UIMzBcSo/K1wUmG/AGXUjnvGMcYva4k4krdebFdFNXO0EqAYgQUMXA1qb/1Nsj
Uga/S1obhiip38pyN1T4NWC3IM4zg2QXNnDkWuW+RpdbpIRUZY1bAFhd3jglBGluucUJ0z5BpM8t
GxvW+OCywcCI7sOHNiLyh5c0BY6Z/ZQHdmh+1/w6LdNMV73BEMqECtGWx1dZSNTvopDx6Oxl1Hmy
QPm8kyVxe/GxAOgFmvsUDQ4EeiDTI09wgPCvw2HP29WD5R5bjNo1d1T78wjMjM5uT1AuqC851Q/u
tK/BSx5bYIlV9LtUhU1HtQspBkNjq6EgWgsnXfh4P7TKxKFHmqGW78KMmovAm4X5tB9gSu2FZ5Zd
BfYYtIQCvwxVoWmPgJvpgIABm8usbaorWqCsITsKfvgrZIyjyqSmcarYNDqQcGsR0eyLEoOXIwZJ
TzrGO4F8hcuoRKa1j56CNcIMuo7XyuMRNQQw5quEfBbqYhKTgpujUHhat5RC4a1UFFyhearZpVs/
hLmyp8uySD5KY9C7JnydkxTbMFquYXkosDZY2rA2Sc7idt0A6RxJ8hGSSfJUbVCetdNt0Z/6whCV
hAtvOqVyz6zsU9+q9GwtOyIKGp5FoFAK7/Kh7E/NM09s0DKiz8NQlunj4eplVISxoMnax+XvgHhj
2NdHkfR0Zf8xi/SYF99Ky+icXzlOgjWr86alH/KzAg09sqAqd7VKAozD6+4yloMUFpKJE2VZHiG6
Bp2nag6LZNWkh7/v4uqALFZ0FMAFjwf+Tmu5QtOYjMuLfPu8CogECJoUbpvQrGi5ye2LguP4FqZi
XBK9Vwx78j4Q1yWYoImODN8hi4zof++SgEdC9SPb4mYNfJ2PDVupnTxHN0md1kC4a9523qP0Fw+b
S5eizNWKiN4PcX1kCMf/7arXRDd2NFyG8CRbeRVSRgg8Z6V0gxY9LeClw0U8VKwNtIRo22R8X1U6
NM/xWitbAreNz2OxKywx9DFyZTjk7MzUEI98NI2myf18+esq5yMlxra8xH0OtSca55p4XHzTTkr1
qk3JDTqfZwqs62nRFb99fn1jIRrsGiII5DKNyF8Arst8pQyxL9mYvFTWMZfi5acrhcgOx74iaq33
Ye0X7u/o0pQKE+kzg32Bdl5V+hlePD7vmUoKjEjA1AujgiZekCzJWNpGrWMTmVF/OceM8O3J376U
xfIjmZLfleqGc2OUcDVrokpNztJ2njlkr0dgaJ4NIBsU6rnyzL6cdIyNUTqjmZrycnjN5C8dKFOv
q5nTfS4480hxTQ9l571Ssjml/dPuidmb8HnuzjpnB/L2Lq/aG6owmTtltg3cyh8elraaCweCesav
3eKaR7cjLW6PWwrmFtlI7uJqpEXoehNXuCti06fu7x5QGbtrRuRMWLAu4SE4kK8P0N7mnG8pxlKC
hsn8T4a02h8BRp58N1xhxHKKouw0ccK2rHtiaMQJCGkH+l04/2onN6sTRimyGne5jgLHrRS0ZAU3
Uv2FUxmaRw6FN6qdh2j79rNEbrx143Y/mBXWdkImFT1yTzoN4PdSjIqoejt8yHOtuhm4H6ERvDj5
d94+EEQnN/Mhj8syaM/RQ6SxANqO1pN4yA09ALuHvOx+WsWiZeem0xIWsTQnzVXVh69AsM6CKmO9
dIZAgWW6L0ZXGkREFDIbIeicWzhSaddAF/x7Mgg255i+nJBfSxKhUpnKgUH3rizvXXVAXQYovQo4
F2sFEiXYG5+0qFLWQ9BxY3/ETlgig0OgRZ0V+r/VJcofSXBfuMK/y6f5kDYsg+BXUqsXub+30unR
kxjlq0dLOyNhDXOrJeaCa0wqivFs+GrYkWWI3N94EzqzMX5AnYIa9REzZTSSKoj0nH3OKI0iUfrm
J31JKvs00sayFRRYLf3oeT9WtOZpgG1tD1fjC6g9uZV2PuT8HJtqC6K41sqgzBg3jw/t1FxGlkFi
cEgaq75czvMjsXrPvxlLshiDMP+12oIWDz9WcBWpZmH0DIznCiTqBYCQXmEYsA5EyVZ4htrFkmLQ
wtK3tgv3SIYsHh0AlXOW9/N0ii4BAX9xKztqlgj4tWx+KA9j5PfU42gCk9tsZ/A48HKHC5m+/J03
+CQEUN2NB2HpMNBRWOFQonOOc+qKXkvgm8PisosC+NUc52ELhvl1ihpc14aKtk5pOmQhwxlCu4B7
CIlt2ztRkx8iI4JvEmRqlC4lSV3bRC9XztFAK8TSoPLmf1ozh58EnmS8LvARuX+O8yi03eVA07hp
D6WVC4BSpNWoisIj52rPfjN3OoCpB36NpUk8ydokcnd22E3KTN5Tx/+BICExFM6NYU5/WH50s2tv
FjoDVeX5d+f5PN+x/dbwX0kveMA2Ga/IX3zEiwYHo/z5XRigjXDSnmqfWjdJT+Y7BFbDCz/y9ekW
LyiXEGWDFIJql7I0Golu2aFcrLauagxqvU26GW0KsiYQ+nntY4JgHB3HgNtvWofFTS4qch4NBmVV
kkPhD06QsKMpLZXePBAmLJfxn7NEh6l/rmq7Seau4YXwA6AvYbB9aBDWlIUaki2AQ2PU9dI+bCNe
Gqa6SAX4K5h97/PQMVTxparus1cm65PUodlwDtyUP1u3u8hUHtlEttCEcQpuCS6HWjciDxneEo4J
y8Ighh5Z4mFCELmHzJKdHMp8jNsxH04HpcuK0kdT7Qn6xsQlr7/w630NszCayXdHX3+HxAyx6UbK
GOo5jfGYWNx+elTGbfLYKA4ojJm+cc+59BHvg34cQ0SBYEILXrIliagS0lF6e1tLijQWj5S+YBcb
UKZN5U0SGRje3Zt40OpY55kN/HTO8tVs6hi5OKSkK5cOGfIVsuVgvdyoWVjhyliAd3Nm2And45Qj
OTwIYYygCxTauIgwfYC1lKA9CGDCa/W/f/4/nTIajYvgMode5YWX/S+1KauaueODAmUImBJXa6OK
wX/Q/WgRw5iPUEBBTtIGXEnp6INM6HBC/bD9qetFG0v+zBhT/Fy7p91t855KlLtUh5puinkwHvKG
Ljsuoh7yljyYA3KQul011BalETE1FRZeVRIMnQ+LWPWBREhn09hZJelqj4+ZWOgsoyZuRbj0aTNe
fOcQ8JCdPAgN5It0S6lnWUKoIM/grIk4K7PRz+S0AssrnLlPFw+fHA9ryiEXHLz/rNi2tail2YdZ
cqX+YD9nIxyl/q4ZBwpYeDAgPvBdBLn0uOabn9wEXCcmpCGHXfY9Z7F8fXYKlHOAnJD+XepnTSyR
86MSVpaqU0CgvzsXX9YheGHyKXsdZlDNPb6njdtItE1qmvw/aFQYJ1FcUwuW5LEpasZ63qLpw0gV
YyOiFpJtPnD7saCda7T89YUw0bPn6EAgoxqjFX32ChQFOPnbDcbk7Yv7A/2VNJ7ZnH8Ygb7L8usJ
jLZggRgw2BL8RPjjIdiDhCXsvtN3DKcMk4PPGPr/0UrTMnA0hgObMzLSYzgzdhpiDe/whKbqZSWa
H6NIWV2c2DxubJYrmXcBlaBeKSWCMDHwVlbc0Ob6/xB7j9TUuXr0+VO0VjWMdUSc8hSBHrwQ1/k2
lB6VHxopnxXuxrAyoSrMAEZnCtjGAtG917RNS0v8Bl+XlOpcEBOu2WbRvapSS/K2iQf6u56omaUN
XkP+PrhzLHDhKXlDdKr7ZwbNFcdQWk/SO+hL+FtVhKTCenkcIfzZ6ZHRI9gsu0UuW2SwiZ6Ir2e+
Xq+jnLs+18/dhefLp9gGOvMbimlJ4FjBLenkCEuV0jLYSKFPRjFf6W2QZpoyd7XHMvCgDIcviWXt
3rBGIVIK2icQbKwU4v0zkFSrEJtYrBJz5T30mb6KwPO5QendphVAV3PDtoeHYYuE3mY4xECmociv
f9U1pPkZ9aXiGvatRRtvdO9a6KriqbaXEP+r9iZDbk3YiXYe/b75JX1tcmIlHosnmNG5d8VCBBwW
u0wbFy/7VjV4jLHcGaLjxRnIbI9lC1WPwKOyQoGXIufr8qaGXwIKRYXuw7O6dmZuR2ae3X5+wfpQ
WxANNt9oHtx8RxfNmnF4+jSb1uJhlncvyNRFYgPHyT1+pngsOtPivFgbsZ5ary6JdqAob7qIfheq
IiqjwA0RIb+c6WG/VWD2QD+V0NDIA1sQdzeVUP15wkL/VJ6oP47/x90CamJdF+h5WBnCUscfAATE
qNBFRb/ZHwg7OllfH6BLiaracCaZX1z8/QyrbGZkDy7x1/LmzJyGl6aoykWkpBvySY2AissCl6cN
CAGkj7w31mL+oudRjPD+R2aEVSk+AyEndDw59+d4totG0bOQV8o83hpf/l5/nMqEAp537+/xaL7s
QzVtRdfPR1sR3dOc9GHXuncnZG32NgLRw7y4jsK9GbvPtlHwPj8S33oEyzMwFS4eylNqPWQmmWs/
8xDMGUD6lvn6mSmyio9RYiLiihD93JClrck7Jtnf4bCMOaPC3Whit6X83Ls5nXSobjVeuIUA8To/
LVkrLPHZf8fdiTe5o8g8dltUAl9I8W4Bl+nyBU60JWWfdhIt8MuTqhd1GABXKNB23ooCVwgd/BqE
3C25mHloRloLRnXsXXDo77V0e8fb9cDLGSY1uCo2MfkQSCJcz7FGbGjGlw6f8Sq6RDUXRdzKag87
diZ/avXPZ+JoorzjhFuTPS512cXfTPnRaG+bCggTJQ2NMc3MQ4kL95vRMWn5BdEELks4brOlbDNQ
lQ9PkI29WOyrrPDaZFogs5LzqThQLLch4LVvWHqBEts1yuRJGH7Ks4k3wGPGQihsCuK7VIWnowGu
95WqTHIZX0YOjFqQzN3cmF4/QHoEpMeVjnEXkNYC1Qacmix3cYF+sSCjwDZ7xlapVh8x9PaDwN9L
yDB3ZijLiDM2kawC1qlk1AH/8jCglQls9lSyH8CuMcoieH/tekT5vk0UpJYi/NspmaWCNmIvUwfO
gM9AHvlLJutecWeWDdOsnpQyB9+dzIwEgA5Rkq6xXWvIYP1NGCkmulX8vRTsw4A/9prlKfqV2JTG
n4YCog+w5mcNmPruwlazeDqBN0DlRLzn+RyHESFIJdTug3pWosGQXs6ppGznsbLT9hZ0U/HH/n1O
dyRI0FNhPzQYGqP3zoy3P80lLU4NiXxP2pCmhq4PicbGjmaDwA+h6mdgYxs4xFmO7xP7sOgSdGTH
Pn4SVTZFD8CyqThhsTT03O8A5WqXRa+9ScJGp9jGExHYh9sYcpS5JB4g55Cc475pmT8mlyXVM3uY
HIS8KZgnbLI8x8RKl178erFNu8MuHx1lO0+pUZ3rD/TsPXUKQ8I97JXDAylYkK2lXczUWBJvWv7E
A5ugj3+RgsrWDZIty+CBSHAyGg5hqKwdh49tlesAzRNM1w3MBpe8jGs7KLqqQnEbIZbJp9ISbSPg
37aAoWpAFkumh4uHGJHv8PiYZRdg1GQLHv7Z67GiJsxttsMOMcfM1ZsMbZzcgZwvuv0gUf+YdWxY
ufSROW8KUGUlplRySYFWeKdAKdi36HB9xvcNrvvVSaO30QNCiO+arRoDYH0lJDGcU9FikAAK2XCb
evcwKijiI67TDE5F0fERRvH6QUChVONBO/NUFWyRrfkEKdvOXReBF7Q6l/zuDfLKd9yDwXIZ/ErX
9VXktTPFsfhbtAz5+7yVoCzdDhSG/aq/eyTwowzEpDoQ0RH8QeEPRlerQNBIbl6TEC4DDoUtFG79
51bKlwzoGPsO1te+Qqpexn0wrUIMk036iRYq9HyHz5eZgHISttKE3VjMkv4ZKyhkyyKT2PAKst/7
aNchny0DmbPy4KdXCBPe1VL2fIhsVCEXAKg0n9CuVhns47Zj/9vTRht8D6jdEb4Huziu3CFxXpAg
V0uHOOCxtZAP/Iu7WCdKuY4UAyL2XWeB0AipzRxPMy2ZIrgqq1GmG6upwuXztNBI3IWE+pM4jJrP
nNiPyRpEh1yFFc18WtJTvwolqWbvakbUhcvAq5uIgYwW/d4CXcOrRgE+jGq3jE7B1cMqfnDlSm1Z
OQbeWxZb/7UcFtXs+QqwEyTIJZa/JBBE/AGEbp4CpMxluj4NAJJk53fhR8YhIZHdO4XYFPw6sF3j
dNW8ZXPAZrDzpGzKxeorOTPtw8iqHUd4S8k+YuOcoRkilcr5hCNdK3hPGAAxi3oalEb5Zv5UgfWI
3nijVrs1IEGmkAKTtxtlNutjFauGVn/sL3BkLTLknrupvritWiozzv3TM/2B/GdTVji/gu9OpUdi
YS6rO4X0M/96SrWhVgvngxIC0eX/ZpoEGYy1CUrvdU3EIC8+I4RYBIzm9o8syVdsOgpPpkLNhV0g
rYWSLW3Uc3OzgjKAsVG3rov8CztogHXPzQL+vNQFeXSPFAnEy4URr5TVcY4HlUtbjtNOobGpymZj
u0ZmBzcZ2zPcQrhM2BLmX4wiVV8nbXt3GaQ0PK7+WXvT4FqOK5ffGtd6d/3xBmiK1eSbzd0VWRqt
bXeG283qBHeXmCHNzve37xQSFeAILF2ruTHkBMbP3UqbQ0lj9eglW33geqVjdCxmGO2dK2E5kx9i
oylCiwLwh72RYznjiTUD9DmWi5axR6wamNMJLCjxYnG6kxGWLSHyUFUJxVItSYiXAA7J8KmLvG/q
zqDszDqonkJuJezA59BKviprt0cg1TNqgh2LXTFoc1cazHnCDdpVT9TKfchZ0cqdwh59zLs0/+E3
4FINnZ1llU52zsPH0p3ENQJ8I7f8aqkP/NkV2QysLms0oNJL4SAIfRLkRBIFbpsCXixH/RF/id9p
InEC1sUsftsC8oYcTzE8uxmEFLNgMoMWGG953aHRb79ZmfKdPebXIX9DxC3fBHtilRtTq1+w14DY
Am+u9zHMKZQ7S4eA6Zj4J4zoT2ZV9PRSHX1FkpJBj374OtEARiDfyW/ZZcVOO6V+gAIk1QYArd2i
xzjLNmH3SDxkNtQ3oI25hrsxMPrKAO4qlc64/Ogz0x6GBPjTeuo7dwfVEYxSlETvI3y58WlmkteK
OmeYkZ2tkVnKos4FdH6tuH/IOTS0DR8TVt/sgHfeYBbtxZ9X2OqxmlZR92VlJmsxvzL98vfXmYza
nLW2iGd2v3ZwRy6cLUYN9uzkuyiMEkveBkG/JtN1ttAXMKQ1stZzPK210Xo1zugaP/ebNMrPWAx4
eaH7XzEEqYI2BJeHEMxcQuu7gov93LCyqbP9+a81koxZXE7OWkFqodJEEZMLw6JOobhZzPiGatMm
7M0X7KzC7xnpoZz7y3ddHbtpaUozMYIqGjRG0ZziDhGYnkN6Enx+mtLJGgt2LYu1quG5idCUu+D+
pqvuNVld/LBNa9HXLVw74w973X3Z9W2b2eecRhwOdWhNwtPx1R/NRF3nKi9kPt3QOHhfxBLfApnQ
zOU5SCFS3KTWlMdQTg69Tp0Gqt9Qq46D8EpNoRxi4CJmz0iJY9qbVUXVLW6Jil+GXWK/apitAsDj
PLKVVTZOQsDTRnf9Hvix0/KgOv4jb8VapUkpAfVaoX1r/+jyFWO5KsRgMYaNdLX48wsaEPDYJa5N
E5Ckg/CL4sit86a39IzApo2u1G/tOCUgp/jDfS8+6hqbdxTejQwKUyIq0vun/1NllVexhHBwquac
l8DG2arkZZHcQ3KzYFBkD5IOc5rO0zb1ayyeJDUkQDneInAfr9Ztr3cx3S2WF+ZI7MZE+UmqPljZ
hn3tkAKs807/Y4c8pnwZ8OEQKOCmnDshwc9k20+f6Iz6+Y5GkQA2hwyFwIIXE6aG1y0DE2xFAJTG
LPKaSuY0GYH49QonpTerZ0kc7G7pNnRrgv++xkr4WK9xPDpISiJ0JL9cAyE++Ta2ZByuA4t9cPPu
kN2+lOg/8hONi+3PL6eLIZp5ryhv+KisE4pI8TvDltLytr/EpRXADK0XOp98lZypm9JLtslwwQuW
B4bnw6irnjDCVZT3BRiNAkpsLBKWW8mCobfFIX+yMTfOoKpBY2fwo7IgG+OisR8K+GKH6yOgkYUD
NVLRvhqRg+VGonJ0nMkvJUTy0wtj4yYGQM/m65sibf3QXZnt//0IVZUoiPkWq1mWNr5sk+7bA/fu
rzbc61Urvl1dX9T4mabqYqCF1olM8IKKGsaOZwAlb+sF5NOznF0nlDhize90o0apnpizQ8gB8WkP
M0Luyeq1p9EmNxj4+uztW+qGbJBrKA+vGkE4E5Ixb+7XkLsXXbrBQBplXnPNnf5kxHBn6LoiC1OH
sQlTgnzTubCnoiWUGcvaFiSS0GxEnBF+SslAj1JV/X1UTdUWNolIibi0LXuBaL2smEA/B4Cfxf7q
b00ianwGBkrphZve947ixLPEbGA1yj7e0JvPMY/MUqCZA4c68+5R/rAaAMMu2biHrBup/E3S+GF1
gUdCHnevSk30BAwfIrjfw3cQRyz6kTBfH32b7VO8MO3Bys+ipsjlFrRsrlCWxpFYxaYReUbgCAUq
5kuccoONCz7sHGjz/x0tiR+ku5scw7DVDllTaKp9tyHhtSIQ7tjPpH2yZJykGLUw6YshVqMYAZ34
s+XNiaiWpai1l/G+1aPQI0C0C+FpFD7dYkCOwVjGTayGdO173TLdbxOYdKUz+AimeJhbeItHNm/7
NgqNQbnL8riy2+xncND8jwgzNBNUcIJBunzsK1qzBwwwyEyjDn7t6ekZmmWHBN2t/gbe1RNxWDWs
yuaM4Lr4cCLFaCL0K09gesMR37dXfPyJTXSBwCqCqjgoLXW3QiaKI8mLAEd0GJanQY/8ZG2+T8To
wOM7ROHzLAZu4o4lMVMDxvUHDJaumYBdwHAPq2hq1S9M/bhV+HyOHJif+I/tBLYaPURqNbxmcqQA
h9ES7pqhwQ4m/lpIhXrB4kNEMfeHzT7JjdOrj+k0VDLAfuxsnOt/zxQYSW1GgHNobs787nFABn+G
Jqh84fW+lOaxm+9uExxsci3O8zXgugdsNIwWrA3YXGXIaP0V8m2JNTTG2JW/LEQ3cYkn/zdOETEJ
vTmMa4xfTmEChl2xIihHQjadD9GLERDLoX88RU76pwQQX5wEorc7BsaMAmXJfX4UnZk/xRDDvoVx
2ax3Sgt9Z7QNqdXCw+GLa8TsraQX/2KSno6ZWsbhPtjEc7eF7Y4OJxCa4U/UBmJkAz3XzpWYped5
MuRSrw+HroWUwHLjOoCNWIPObIdXj35FEffbc4cnOZuhQdh/L5tf7px4RewCvIh6qpPO/2TJ33Ag
VESOgBFd1kzaw7iNRQ1R6EXJ70JgXTa3Hu1wfdB+KzoYLTxNDNbXZugtnDB2LXOB9Jx+UPjfva5u
sIsw2Qywx+EcTh0D4+QhNcyoHJBZtf5Hrt5VGkun9/PprgU4JJuao3MG1LLqj9bPP+VnY0E+EVFu
sJkujUr/Tefn4vZXsMqPrHuAz4G4h4j8HmuqYLrVbK9Xv+wuchU3+QBx8ABqPfBtDWNWc0UTkc2z
uqkx+xD4rKbLH1xHPZPZtljcBXTiA8PgrY4QzhZQnth4nokXlo8yPJwPHlNwt4CLl3LW/W546QyL
jCVISBJdSwIaAccX6l0JDV8fAuixvrGN+nmwvlVFziG0dm3IspPpC1sBJLvT5lcgVw+IvfM6eTYd
LW3jPaSWi4OzX99WJecbGa4yq5+dmlXx4u9MAboVDd8qERfRmgXTYBnD27UQPxllNnrlfbtR+YGf
/1qgBvotT/4NhRuQ9oanmVzi9fdagybknapBpr7oP+drit3lCT3euqzZx9dqVIEpFIcGY7tfigAm
S3AvFap5Un/MWKcdkwCEk/Jak+DvJAJITl0p/nl1KVoK/M8rDF8bfDVObBz9RMKNJbEzEFHJs0ss
vwGXWgI3Gc0EfApn6iSvQTVumVLbRTm10Pdh7KJ4qOjonNdRDMYqBihEp2/9Ne8lN9MS3dd4A8E5
mVonoRau69NeLevs5zv5bB4ABG3bSMTzhDMVlaU+SOYwbHvonZGaBGjVu0AAcpZWdpSuGwpBpCM8
YwWadFFaRXqdo/Os7LUfuKz3sxnWP41QG3VMotZ6UZ+H2+AyGnplosaMxEPDZxWY2yXk/Q37jqr7
DLaWAnb/GU5wikJc+wA07joR88b8Gjmn75FGiD4aP5MuzbXOW3mktjNoA/i7GG1qtKtfpA5xbWEM
gcYwy9w0v+lVvTR3e9B9UsSH1tBKeU4ktmatOwyDRat0u9n/dH1ZGfzeeC/BtwMM27VzFWV8n+8P
2GSe0WSCYla3wUNuVz/nCyXY87UGzrBU5ORIQfSjourKofEWaaHBZpLWKVGnD7bP/lCoditrP8zd
vGLspv5Oq4aRioyT4cxq/JrD4w1+XlGeHM5sRq/QIfNmpppD8Q6th+nG9kU4iZ5P8SlVqfch7hmR
FxzFRs9TzukKGIKKimAJwc7b4h+IKyzgQLSJN03ysS+Me8GKHuGTHFVYacxtNzTgTqTAtc+IyhGB
XNK7X71Yz4PO8UixEgxI2o3n2cX3AUXpKEBewmwITlt8Q4W9mrljdZaGasSA8w7tspibOWGFthLk
8beK1sfXZ/5RRLkVgpi+qaL3pbbF13JDFGp42lpkdcAy9krc6akxGl7m/WSy+csp93bEWjqYOCCH
Y3fLLc17hXxeuRDjpJpZiU1IcUgVHkSczZE+enMUxklc576yv3KsuZZ1eUq+L2hVkL0uhhbwBQyK
EgkBjeQAFojVjSSa1sQHPWXggH763nfdBD7N3aBODkNuZAhI1UwMp2EqNa2EiF4Yd3Dt8ud4i97G
t9WkLU02gKkuelwjN96cLY+fyPpMraTwdJZQr6ZaB+egGSX5lwnGTaE2v3rWkwkP/SSdVqE31+IL
QajenKMW2/3gv0YPHBCASmi2aly4P9SJED9XzZDewc768ku6PizSr9pncQvbEIPkWMsnhAst+XGW
F2e+QADuXOlKgUHwWboQAjfynI5hWVPyU3fysBHtUyD1TuLZ1e8xe1S2hTy2+Pux8PaU97GJjlzU
kXJYKkGZi9N12NOv4PsizbdCQNifef4y3hFtMuEA1EjM/UQT+TXTFf+XOh2VGs8GssQMjc7nzl2L
UfGifxJJFG5fGJRO1NMia53CxPMZlmgE16HCpjvwxnVeTruCfFwujnN1EQmI3rDKKhDfF5qRITNW
1eoGyebch0qX3Lhv8ssmvLQUiGNiR7AmM6PIgKdX3H66lU4N35Mq930+C/UqugQVoENSCf1NvZWu
LlkBmDQjxj0kjecf90a8y7+jwnF6JIf1dtgLd3FqAmOaT62vh+345ANfwovlI5ZXviccle5nJI3c
xG4unwj/1oqqlKE1r/zFMMlDuT5hwCGexprg2LfpS/nWNvuA8IwfoOelb8aOLOZ5EuDBBPMFT3qM
Vyp/7uUKebikz33pPr952cqmVVNbiaghquw7lehlMT0lDOdk/sXMNZO5D4+cStWfgngpktNxOHTX
KoPt7cDTN3mSEJVV3Y4X6TrGk6ahrgNlLmuK6Ymagernj/PEQU0YVKPZ6Q/8Vbply3vCXhyO7kIY
qgNpbRTaNYhrAOc+M9UPYGJ+mgdu9MWjZ0psAL6BH1CCNbe6KnNe2d8P+aZIQGSXpdoPphmvnDzt
ElcZsTUOqDfeHGUW7Gjt9beyZJVAkk+bMQDfGRZ+naJ5Mod9FYN1lRSTaWsKouM6m/h40qTSYXPP
0Mt64HwI6VU1XgzaBwVJy5k4D7ANJQhPRLwJTJbLtTeTZzlVnzzVDbengEhYLhb97tmfi46u6bbv
CuRMxOgQ0VGXCozhPN7WiE0llBEzWUYpt9gVAG08GEvxCyXATrBzWaq997SaU272LaTRCdxZ3v8X
mn1OJLPNtE63IxjvSjHedJ7ArSsj51Gk9VCfiuSbRaCii2R/lVWelxf09d1prYKhlFKfBWblTw4c
jePUB9JJE4x26wksgsiF27WeTe+ooI4LfsQvV/yHy4jhkTdkr9TMVtVUivehkPyaq62dP3Gf9fIe
KEl4Y8GNL6EKPCA5R9qzJPJw8FQ9wJFBv358XuPH9hCFiIC7vkWoxQ/DruJMZei2gpSqzYgrFMwH
2Jg8RdYgqjyYsxBvWfjbFr8Qn6z/72RxQUGYeOsJ8LJDl+JlNrGCXDQFTePjyDGU3BHprZpEX7V6
Pw7Jy9p+A01gOptuAeVfmY0ss1nrKeh2/9+HnfjlupUl4OFXMphJx2ODTDxSyryaHeY0e60MuvRo
ShyWF3ly8YxqVOdWif2hOpNGBdFSWlqR2+5WSfXic5jGmkB6/FgcjS7+GXoxXIFTGDOdloT5jhd2
FCsJTXSNT5jFDzY6j/DmfwpkDLKj4olXSiwr2f22vJfEr4gd3hylLAGGfACAzXVsUAWanUA11gg3
92fJS/XgG9ebhgSJfuH9fvEaTYWPWfcSTLYB1GFNCRW6VS+X4/PWbvlXt/gzyAe5jq+LQopy0L4F
W62z3EjUQ8jijPh9oJrqfndCEsMK3YSFDyxKQI1dcPwWV97sCk20Ufqh8Z8GCoP2mUsTbi5W5a01
hhKJqghNfE3ta6gGkbEupaW9sLu6b1mr+HZVy1ciQTrkx0lTN9krfg+a8GLH8hAWdstlkcciYJES
6SnQbZ8+PSoHFXMuFUkk2jlzUBl3QPBgqQz5+wKtzrS+Wn1IfxCPUl/HBPHOMFtErW/0hl9XzAVY
3BCRRy3nmFAfTgjUthZgcl/M6wbyN6BSWJI+U5O8JpwzQrfMT+SHuyMjZ56Tv1/ARJ3kbRYi90Y4
kKzS5FjTum8iXblzhjnxQNUzv7NIAr5eypKKCNcwlvRRii4xZekoxiR4zoXKvDmCMOJDtzjymNuB
q1EnOz2q5y5+4mo1uXH53ACDbQKoXei8XY0OacrG/mKoqKFYh8Zqlz2uuzpORor4u7iFCsdyEl7h
AqZgOClFjAYNUliZd1GdhGNwyeD1PommpzJ7vA6y7nXjH4a7Ufk28hJsUj7m+aJsj2yCu56V0dgQ
xoLSfdN14Q7l2uMG1lZiZHVyMaAkY6mv8zfyWAqaYesMxBsArOQ4UJGkaQzyP3mIW9rXYXvBVKEL
KLBKr4fn8Vrl2eW2koUvOZH4OKV88xYxJNp1PqyNk4qSgaQfinSWhEbQsou7sCdbfkSmZsdy2lOF
hTbb+LjitWrqhroczybNHO0Hu9IDwdzzWcjtrt4iBrQsv2YE9ETI+/ba0Rq/xS/2a514cXjvlLS6
FcKRG9xbMycK2jXmRxx++PGwS22kjYyhltXesRQ5FfzkPpJ7vV/Nagutfw0UVqsF8yZ1aczEmVTH
4sq7E3a3l+ppurtB5gbPH4aIMVVBkuZClpju6r4c0WCxf7X1b13KaOHaaNuMDxk42cDBzgT0ICap
sanrEnTusR17lnwOjLffyKuFSQMPWIVzK/xUPDD/3qiStuWsdU9Qb0v6GhvvPd9Lg4SeizQKbvbx
q4vIE79jwlA9gHKjAhxlE8wL++K5bqr7RBw985hwvfe1nsV/fm5qGPF1G9yxAZvJ3W/uePmLPwUJ
Dvlsp0rCknExExDGrkv4SQxqlgLNfuDe1m+liHb1Hgkrzjn1uO6n1ciovnBDPn7za+VKfsBF1HnC
XbVXLQGd7o/tRIjcjKsPjhwxHTtb6gbSYAO/TeC5cGVbjZnNheys3TwHEXyC0sYY202GPTwzeabQ
IYBaNDQgIT6uK0Nj3NTESK91Fgd1I0zAGYNJ+zcIh6uaIqceP9mue6jHZSjtww9upG178ZzgBjyX
lJqZaDjvv+Bgzg5QqZREXOshKJL84T4LtIX8iwv6DwwDumvtsLnD/EBqPRnUITh2mWBbtTLxuzBT
ZpaGNAXRUpnGFsuzSH9TcP0iQqn77rpeFDrj9nA5B/zscIgwR1d33xTDU6jlbx/Q56V7kOyjuC1f
GB6Y34lLWPS3TJSM7+CfeurnZ2lp/Mn9ZYRKKsSUmQ+dHoAC1kCE2lwW4MxI7D57l5jw15wQZHa6
jlek4vLYiDuIuK8X1bv+4f4kmoZw+IsuPcc/AQJSfRQljXfHo43SFuXgBbtHNHEjJu475R55pTM8
igYAfKE2Eu9lAas8tRZcIdn2KLKKg3eG276yED34qCFgw84SklQQQQ7rLS4ZcUh7lZCdYxClEal2
vx83ThDHvnNr9mY5J5zxdBm5hwoGtsKhaXBWf1vX6cq+l51rjfBnvDHBi8+OjNbQzmz7msR94rcS
Pv8+Acil9W/RDSrQ28ezng2u59bpkn5YxWmMe5On8wYYnrFVbTHHfk9udbCkBHtPBveR8uAsDDT4
4KfZAMBm1q2xUMUwMwhBDWwKfsL9X64oGs8SLCuT3+J1w1dU8hjDWx9lhoOkhPVBEw9o+tED77Sx
WD9O2NJpywTQ/tADiIW9vSnPtRNzvFVckP46RnP15I5l7vUSqqqp+3UNsdbrTVTnQCA67O7fUAyN
9vacvO+Dt5hxzW9Fu6btw7GOJuG5nASXnLxlwflprLH+brllDUcbwlAOaFKdg0MVCxQqVLc7dedv
lOZ5sVBEit7ZQRm6WkOzp5n39YzeHyErw6qh0++bt+RXKe+YcWndExKyTKIbSR8O/7skavRGzurJ
6+7NBacJTQc4rSaTiCXOBdth694YObK84zTcgVJwaKISgTl1Oi4/VifjOOLSnwncZ+bSaz6sAGM0
sPFlkOt8LpVtotiePAf7fQ6IV8PtnDA/p4mnGFeII7ab8uv/+VpuddAhnUJHXIlAnOJw2uxYdJQB
zQDBLmda1QkIL10emyxbH8NVRK7jedTcNSk3WXK4OgkBqelk3cr/RcMCOkDNHaXfWgluMo+Cf/tX
i9PY+f1b2K5b0tzTv+X+WAvvNxJ0TDelEG6NhJ+ow6yQ4isZFGv08YCnlxkt/GOpn7V31GZIllyl
DkR+ccutXM+f8QBNUq90YZYDUw/sGth/s7YuyPNGujIEOK87RxiMRIOgyWENKoXXKFFd2Hus9S6m
o3Z/7jvARNVpkoJlYHyMN6j7YIwB1UTrNXJF3efU9i7l7fS11/uqLhAe5oRnjvhE0fuPgrr+2dA6
O+xzOVZrt3iRr7S1HM+4bf/YftfrI36S/31xo5uM31+Fc92L3J15NhUimhgtvUUdiV5wkLHt1rZv
bgYip+C9SSTcuNPIfI7lF7j4ZAO8Y0Xs+1wGxQ2XlM2op/Ka8R0n8C3iAelTDQajaeUoq+OoBYPd
SHSJttnh67U9mX/AX28FNH3Q6/uhTdD7JXLvKiUSEIUtDJDLru9fSI0So1b9Tl4q/zEuSQjUsni9
KQwVm5coFyN8mqVOUCd3q+DD/6sJRfYZRcGwqVfRX2JbR4Zf9Xvd9Kzk76oKWRHnAs2qSwLerhUo
kSOG4YUl0ZI673h6sXIk5XYTLY7yc7iCXZtCAft59yf2fsTMd20R0GiGqLPKajqRuXiNlxHD/tc2
F7p1tKgb37S+AYEKKbkcIdEw8bW/TOUfot6sqIpo7qMXoVKwMXllcqETUi1ihMrA4GfJ6k6eK9Es
NN0qOHXMKEtckUeLhVDKaFJVCj5A1pA/hoHM9V9E38OPbu5/U0MSAZPCoxdh4HdeAMt9wQLMmcNN
/ZTmBBekRWvQe7s+AKgzyj1jyayYDrJglxTmQjeqm/ukabqjyOCylQzQzh+6elQvJWwh98vkcGI2
LnttzM5eTsVa6ZF6XnWpWlaFspO11vg3Ck7iuEGWIPzDl/KaVM3CgtcvRy12M0IxWFdEdRaGQmcf
QgeaOa7o+xX1e1KsSbO3pLKTmyqUXyB2QysO91fjirp2qWqnyDZRBowTzswhU1tW9Lc7HYCSqq4N
Y/SfYpBbMeKq5SUO6IUVhG/Dq2mSBocunLI1/s8U9GnlRy7YSIW8Q2XQheUzl7AkLOxY6Teh9q70
IWoXg/oakPDnbbFOuCqiM10kEK7iQqxlKupiSli6iX8BkSkR+cEHd+iskoRRdzX1VULwv4Vgt1zL
zLV5DbZmoAlQNOT6j4M/A1zAEOmADYJNEldgJC4Wloykmqiesm5fTSpgwgygXDKvlB9YJCg1fovq
SGxtLiZ+IpZPrgFrFOk/gNDl4vXl/SWZQCMwqR/x5mhplSwNr1OnLOdTJrKlzMcRulWqdC80LEyr
Z/1Pn5eTdHa4tFopPS+ygs3uPY+g8xoGCe0IsiGXLASR+BghMR2qUIgDsZWcai2qyAJpN+9X2EQm
sR51c78JJvk0in9j2pNKWkgyNCmNpDfKC6wSFa+cyUBjM2lDErBDzaTlFBnJ9yTaY9EQF+ifDGbB
aI0mdpQeHAIfDU0GJD2/xxOI7Ubw6RvmRqwOyQctrngVeA8+ljqBrDjhKf87IJgC3PBj3bzXp7xN
A6bvb9e2fjjlYzHPWn6fic4TLgI5i97AKhwUxFeCFRGnJfw5hXPYaEjVlkRq4AhdH/wVC5BOTqij
eQnxtjetvuLgfImzsOe9qrAcqB5wUE/cVhN3fWSmug2uJp72gxUDQVb1ay2OrB1BJW/8Fxnglp0q
7PFInkc2tk2LdVUv2MfJ0p+58GJxOFK/Y7leSHF6SonnBg62Suo7UdaCFd9n0r25VyYFXvquY+gG
P/k+d2ETDa/RGuYu9ib9W4nbBGycWL+TM402RxhlWM1sQTUqEthuTXuPVHXsZJa9Uac6Xb0j678a
oWDo2AmtRk1uQVf/eBQbIs7jzOO0J6aPtQungsmtcYxEirnEYJiHrxUeDJ7Twd71+URCxNuY7jB1
XhRU7m5FG8HW0HdbhuIkfY56TVG6dM3GHkJfZtoRAh/SwQmqZbqrmklpz1HHTGiJpb2WgIb7J+Hv
2ANl+PRXuNcf2TsiZuNgumsLNK3Goi8VmPMkJsSch4OPyN24UnUmYKiZEd/P2N92jg0vHmLrEfS5
bNL93cRP1UmmVhH00W6gS1c90xJfq0Pu+8woLgKCshao8co+ZWx3f6sWMOOxc+AJPIxmVYyUvMV5
YXjPr5kxwhz53Asl0R7azpvoORkunI4hQkk/CR01al/a9w9/IlM7mxDP39T+x9dU1XSER5hVvgZF
tJZUZGQDnPL8accZwMP46tO9NGS/BF0wtsEayGWxlIkvDxCk216eKweB2S58GLOByV3ingmfeVvJ
i6BvFDx6lmzQKUB3mHqzU6sd9auv0+5dsB+DFgYdsGwckHaxw3Rpn27riA2JOnO2GAkae517qU1i
7F/L6IneUugL7U00OjW1MlRdf+8Vi8fiCVBkh3VO//q8kBF9kIG6/IjQKH09jWMcetNpzp/QoJdQ
QHR5u+dMYTp6Xf96oBm11VbmZAusj5fpJijMN9R+rdtww70mtwjrQvaiEcComMdEY5odbmqZ2+UG
j3q9mv6/cLaJMe/MTtyVjU/J/X1ibiOkFMusLjQO6P4OM9UnJFNX6kbxfeEUDL0qViFIky+0/CfQ
vV1QsDBE6T9PpPJpbh4uc4YDzkb5JBTzBNCv8IWIIXcfZCYVrOf35q/MdyIXP+oQopAQtfDg1C3E
9ROGvkPAq2E7GTxSFx9/MxI2jFINLbb8y0YI1DbE5MdoZ7h6SNhMKn8G6Sq/FQCGV6/6HkfBivHD
bZWvZTp1qgGvS3scYULDH2WDZwBtzfC2JloY909JpKgBbaxapEXsvWMRxTNImZ+2PUEuPeqTtwb0
t4OwiwtvRdPQYvM4Z3WPcUk7w4uhXYgB5VhI7HWaaXn7Mvj5+Gkf41zZYHoZGj3l1y+26W4PA0hH
WY6+JBrWaTOYhWYsjgiDGYqESKA7QmUvNysr6XR5HMkOnaiHcDetnDQLewYyn3WCPZvjCSvkh57T
NUHg6tFNEf2Z7mzV5Urb8luIlC7Tyd/kZ7ehzzitMdLIrwpavc1odkgHjB80cwvYg7et5Caf1h3+
ozWRi7TyAgjhVef4QacJEd0Daaimw+/FVYtTW2q83aJSPemcDTmG8/JuhLM2SWled1IeU57iuMeg
SD5jQobmi5OQrpqL+PyTFwrmvUGy4mVfxtdHRenQo5kXY5xb0/yj08UsmGpP6t4pnklkZhQ+UWcp
7yD0eHGsi6xanXNZqgOQxdGZztzVeMzLM5bOKCV4C+y/YtL2xlgNwJU3gchaLsHcZU+/CMx0yIRJ
6ypOkykA8LKP0PWDL3Av2wtf1sEueqB3B1Ibc27uK7Jww8l6ifGPGnbcKYwKwXL2qM8sGlFfpvg2
nTTGWKL4bIK3DuLgLrmjV39X70h1ZjJlGzBI71jv4c9Xal855whlD0VLiswXKR8EIDox+j2+sDGu
JTeYWvpsWlpoiqRuKxRTrzBAUCVSN46wRMpXj/zAMjzIZOsADRcfK+Yt4B5bF3cWs3iKv+zDAKdC
6SlxZUz+B0S3+hGicCB+tD9f71gJKBiCt3sRX2NGcDnfcYJHjVOJvIXiDL0P7lqsi/oD3wiLr7L5
coVEXeH/wdOF/9R1meVrTpvZd+jEbD0Xj0kDWPdyRLnVr9k79vmMxTPImuIDS1p7hoY/wPPpivTM
rmsh6VXBSHxIqKHnRmaDQ2ci1dYOiYnW9J8wzleVNcsRv+e9hSVBeR78D2wnlkCeT+2FlNlRvVBr
qgDuqkEHUfqoT3WLC0Qr1oD+qdALCX5e35ThgSIPbWJcUu5U/HZ2cTn09bqvon4BEJLkArlwiZGN
CCLBxvp3fey7LqTI1G9/yp29ZmqRWtk/uHKgIGVT3dyTOwZEZFjyQ0USBm/SktAxUk98cexe3jMJ
l0ULbmzdfi5Eye82Pt53h5jksV5fOCOScNA7Goo9ZGFcZef6wD/RDUnJtAWzXG0gifOgPerSU0Kw
rFocHjkuzsZa5cI0n8aZ8qkK4Iu6VA6qCFmUrZ75PL5T4KxrukVMJengQKxlwkFZmVARxw5qm1jO
Xcyi/o/m1ESuKiY41YVhLgi0OqzdKq4J8teE+J/I75BtlChT58OqZAOw4CjKgTJO3gd0jXZ5CeE0
8oQ7HXfbh50NMqvjX3nfmytoczqz/zYNS3SuvAx0+tvdbvr8rC9MB07bDpibYxdP77NrzbT0tz/y
sy2fpAyz0/FsCiKGbqiIV0NDWbQUGnFzeKvFQr4xUtuIKxddL8G1vKV+NEGIh1xUeVI2rmPLduqr
Opi3bPglRO26JRfShO+tvgBDNJqgMdxiPAXcS9txJCZw/ra01Mp378BAhw/kDfD79vSbKkvI1yM+
ITM2XHnRcA/GcotObNq8T88cGCK+cmA0EwaIwikuhwO23cOXx5aW81lE9Jp88EYsyUccwqMSuR03
TqmRkbcX0rKzqxYtsmrN5LaiNHVpzyITvCicTQV/naSBTOLLKKMKpQHYHbBEwXJ5BWhmg0MKsxLn
6oJSYxOfonpMq2ge22UOFh8GDSGD6iZrG70Rwj0rHqOweL9XFi0ObXc6L2ABatZaXTdTW/l0zrkN
DMiUWi5PdMmQGiGn+wE/PIuid3qDC6jtiyYew7VBgE3oLm/8+ID3SY4mumJEV+LBT5k9KgykRCtW
3Q93kAuvZ4km8dCgnXIO2NnXnExJb3W6DC2YPcSUFPwZkXtticVx4xEHU7oEJsAFLaaBOEjBCJBu
ZOl0G3MOlw/S/xZ4o6JWaOhouEwZ7P6UVgVGqDUhpBXYd+T85iGv3adxZn1MayYa/3ZUjG1hcln+
ZMWwmkuOJzkSQypVhaEkP59Y3BthoTsAGHAKLCbNuvIe5PGSCSuEbNsiruMdwW2ayVR3NjvREGZy
SZXjPLRt85FU4Etm4SVe8FNqu26l6mYmJyzTvekSLzVxJKUAxKXp0zKobdnWe8KmpPrYIK8Ug7F8
31DLq6NTT3SgZCFRIo4dHIzzhiKlNj2SbOrYKcQIVjvIjnAzgtiUnf5QCPpWppicxfVmAhXXorbB
8kUDEO17jV+cFpQoOKosfDyX3TAls5D0CqohDfYuwJXdRN8Vzlv/+FzSPix58cKK3lupm7zWOC+e
TbxkT57BHe49nwurbzzsmdnG/osY+DRlfGZ3dLZtegLAr5FYfAE12SfUgqvnx5abYwKPGhUwhKAX
CyNiZWtq1YP7q7NMWC+QFN0Xi3XDTDikyuci6bQ3XA2+Xg/yz/RCcb/TNDeBX+g+lk8FL4bJNL3c
4tqUIOW9mRrihrU/RJhxykozOs5E/+RlSoA0C+7DDYZcS9Lxc/kTBtipkyK8XVissm0dMbVTbTWk
T8Ye+LRqbrROS1S+RrtAAG/qMfGa/6dQRq2g/oGa1gFs5nzQaEQWjItgz2/SbJfxr0PcPZLSrArH
YWCvTEjFZrZcxwXSK5At5BUhUjLxprGfs1+s7fVrIOhN4LLl9SF/kHQf9Fi8A7/x2DoTYMan3we+
a1gFHtqEvDj66KmsBiJi20sauIRjHhcKiOif+Vqo8PkLRMIRVUu//rq4UP8hfUd+tnNfKupWQmge
TMl1Ep8qrDp8JiXGzr2xoA8Km2QPCvAGsgBYRKE3hviHRuB8tVElWKLzI4mx6LZvBZCE0kx6e2OE
nwz0hYCITG3RQbc+2elgF+A3qXlnRcvmPVrElUY3Fr/S6dX6HZIIqCTX25oICWSENyohLlzwsumX
jLjWm1OSq1SdvU2VJFOCMw/fNGSg9QDhTBmMKrXF2XIKPYvkrqivYkp4zLTN3LTd5nZwNXTjRtpa
3DdrWahLPYh3Yy1hzIqmrED8zXcchMJj+m5khpKFYV5GQxZdlulKhjRCdOEF3VTe2LXvlQNOoyIu
jP3XnSMXRYwl2aCgpmMOYwkCfiAdhiqxTX3GZNu6HsKBDNRfIrjtSd7r2hBBSV6tjJWIc8Zp+p35
EY/TZOMW/TdDyjFH4+XAh0rpiAl4Sede4MddcOGZtsGqUuHMoqK01Ye7htfH5MxkUA5jO91Krq/A
rGvIw5HLjYP4NjZH4uTt4ihNrPe6I0wWCEhriKw3lfKQcpsSLa7DkAwj1lrsDv5HWQUT+qz7ZqFw
fyVm4lOhTbfcH5Z/Pnv7QW+0YWUm0d2vm3XI/kYkoeJbu+f2KHsWQymJFtwCmym/rhA/cMRPHf6o
CAUhIk7SqUlZFxb3PTVJ0yYOTLduOmd6keN8yuZ2u+2chOTnV19Y+sdm/XhTyefvluviYKxL42Dw
pWDe3CJHFSOhpVlsz0QNEAgMtLgt/bioMxFQ8DJHzXXzl6Rl+xoLDeCB9xxV/n7KOBudu+MsxxCB
ua+2YPNgVay+M6+PdvXXbvH1cPQmkIwOaEYOxlCEGNmKxEmQGrvSTvdMbkye/2rQ4/YQu7pYTfwP
9qWXNmufHqxZbnhj+xJ89uBB6N48cF7DMGwQ/8yxqTXUynZuctTbrrEbWQtcTCtUF8FWdZ946jbU
txF26YNAK1UAKhpxiubwvM6+1RlyFdykZmNOSAdcklWH/6al49r60Zv3NAKTYf2fVkAzsaBQkfj5
Q0yz332Bc0h+tnqH/zAQauTlEOAuYjqVkdX2Dsf1A4dGk3Pyy4kZOqUlwORnFtpm950WV2IE9ghu
hlPBC32yoMvyVO0sEK0cRVPx81wCSqyqHiBC4z19o1bmzFVv7e4fvHFGa1f9NAYxWw1JHHWhcTcU
tdlJuHjSBfNesG95Enhmw0gPq8OVaCor2rP/AHjNlyOI82Q5rv+/3w+ryNUlx7SYHVIfTHwA81j8
+kLan1ZGvkgpsbfP4Non+Qp3nQzpkQVDFR3DmetAgmIMk/y0FtUKZRc/d+J36Vphf1V6h8qhKfSO
2/TYQNcjdsuJ1+MQEnf4SRSIJJHLvWwkbdIHG28Lu5hNCEZRgZzZM3tkPSLsIX060zlmQcq6Ev2M
QXA8MvESaPTrtiw5ov6GJr3yNDxT7yV8RSSxiInxVFP7NC5PBBkcjJXIG7LkEzwqIC+O5ka96mPa
xkWmXC5UCbXEZ22j+6po8fa53Bayn6m15O4WuLClUron8RvysJ4PWd0z9GNzng9bzrDRJblechg9
qO2xHAqcnzifrkK/Czncog1hYA0GhSXD28vZj1WYCRBqsKGrck+6t7sBVbLgS9DpQMxazu8llqld
snFx0PBnGYRYvWsB6OYTUavKvSVFVTl03hi7daaxLkzsDqDExBZQm5h1uDSNnqJpLv77JuQcLFfu
YB4KZsssicrk/NLwEKOXspy3ezC74kllO7MCM7T634dKzXymBT6f6a7Jne72c0SUAJr3+qla8zLa
WqTj5zgWS3hrDANqRO6XJfyX2KGBn4owNbrBUvfB6kuStF0o4kQ5gMC1OYrJiQJ5eQJkgKnsXmNh
N6AIm9L75XEWAcu802GRX0Hw1YRukTYZhCTa5ur+mNKW4pl0fHjAzJEJYmVZsvBtYqPQwM+dsT7C
h0tagfacaye25ejC1umZbrmcjUAES1Y0CHlcrtP/+T3FT6K03AKo1fsHKWsxOCx+AoKSLHVFnrca
d3F6WvxpBSVwKRhRvqcdBVmrJNoSUtzzkavCdGqajdYo6b9AVWB3F+3KI9A8Qq34RvH3E4UAT2Ie
ZD0Z3QoLtS1K0TJNA4Kj+7etC1t2PjgVJOjENrt7kJm84YaybvTfXW7ECrnJnTb8JaUc0EsSLMum
bgyyGoGeUmbSif9dGWlA43izbVyxxMe5/H1lyclyCmSYThKlqwUodTmrPWc/wfkFQpPX6HJBW0km
je27MHVPvWUP2CvsbVGUoxjMXk6mA2gAZ/zfCqxY7MnWXFMdqfMwFvsB7zwIwEOr088wO/ritnTz
TjXh/YWhxDfA7lzVdw8P8LQswEtOt6MkDVLsH5HD2J9PsVhtFl/iAbPNiHS9Iiy6HKiaVBopSXGt
tbBqcqMHUZJk80RXyNpMzcAkogqrrXEeQ6b3DSOqEpnEq2kI7R7rRF1+hdMwZGqXeO6FjCEFdpfT
/Ihuvv4BMnBvD7N056WlmKP/hG+qL0BzVVAKEjwohATAi3eyhKEBBR8A1DVZ3eDNGZNlvf/cSGqT
6JBdVChZnZuFP0t7qw9cO/5xKX2rV1fIdu8SKTVaKieLmpc6e+zhDFFqE7gfNIKCP0vfKWlgp6h8
EG1go+pf+t7jq73GfiNg09eS7hqepyHdnUUwepAYB+1GHgi3W5W6zUr1yHL9MQaXOnSwZqpUiUp0
T9CVNnZ1aCbyPecXGquJbqiOYot1ZXia9jfMEEJQRL2wQbwoWC0aRbdI9z0oAoi0NJIEukyuBpMC
oO7hkJRZaIbg9rSJDpAqdDisVyPsQlltsWSVrNC8WMC6yNkD/NxPsTulgjgXdezWPzvyMo5QIC5m
4fE0819os7xdF98dJj45bHacTNk+PUvwDl2Yk328K+0ZvKTXw1EUMoU6KM1y56xYrS3JBUXnqVs4
A1vohvi/FoL3QZys2AGg7yMrkTJU+X4TTl4sRHCfZXlBkiTOQYqYIIN6PnahLxQkOVpVyk/9Xh5w
hLrb32rw56wCVbY/iIgATBySQ3d36DdPS5iYe5/bKeur7GjWQdzD8x7jXDD08Akbz2EkOn9HMOig
h6BUNNW1C66h9nb75dOhM1rmQIlMnf1m7smHOWiB4ybYeZK37XrwqLTeSbCQHouXzftCmQlYvjKF
mFBI+ognLxDRFXhhE0DoZmWvrus0XWeWT4wMa+ylWiVV/bt8f85pMMWYFLot8p5cP7D4/wAAuoVZ
DosCB80V7j2VXngHjxQYuhAd9xeGI6WYYtfja8drppg6AUUr9PLCu35UUkwuChu/Q2CHrZVc120A
qXLy8c3+VZhdzEuxbv6ZZQLYZ8nJKWpN4fGHXYSbalCprF7/euqzJ4ypdqbl1T3pRSRQiJ/4MjFX
n0OdBBiZl7gMQHifR6ZSW+s6CrJevLg2yBntaTJX+uOQvxXhPGrAdV4q93WxpqhIlVDuFqHLrMW8
ociHoQ1qwgoO0tPhwoTvgD0BlRthhJse4jjRs8lEwQqQoymYvCTZIso1+5hvW8VZBrRrBAPCaY1v
vyd8Vo52TIe0s+x5UG5vV44TLbEwYgGGCaSSnSt3awrxPiqwlT7iGlL+j68sPWwo12g/1yS9/1iX
kRem1Lz750yKHb6AtnqUZbrtEyfLMIjD1XQ1Rwl6k5t0Q5MAtbYPLzZ5ArGZeTAcSQC7Fbx/Tqqi
H4ok5nlSqWS69OJBFF4jDFreSMmSTG4sy2RaaeVn3TWDPyT2X9dzFM7W5mFytr9ktWOJ/Z/LyM5V
kqysQgTAEKdDFC7Gt10QQsOQiMWw+kUd4geDirRPvgizxrX59ztayoOBNlXfOLgqb0ArZ0B0Vb+2
RHndeV1vjcQ/x+VvVtnI8ze/4vd0kDlAt4dVsLUv5wEveHIi4uuE1C5yDVw+vkCAcR79Kb+nO+o9
okQIGll1wvUOduP9Q64fK3pUwvi3l9HVAswAnDWPglFf2xZEqEh7b/mUqvhp6V7hgBZs/BkIa0O0
XdQ3kwzE24X7g2IqBtABmZSa1S0Zg5PImzhYfQdTR0qZqxHeHwKTayyr9Q7zSZx6Vi5yAaceCNp8
2sDgwtuUyIeEkaVIFlWFBOnQq333Jh6i31LOVa6WoVx+W8RpYQjF5iplAbkR6YeHkPIA2X79WWTZ
ACLnHGwbbvdx5FtsZgg7kJhTVxaLntjdZF7eHAvVSLr1GxSolaEpj5F4FX0cNs3FXnTTEy7zKf5t
o81zVq3BOmdEm/mayc3goVCJRhrAc452F5CulAG13BkoDf7gyNKB5RHwiE1GpNQdAP3D2jB1Z4+Y
8AKxM5a3T3JFCVtLyXTtVGs+arZfT/zO3SKfnPe/B/97sFnPNaPMiqoyFg5OaDH7OApiHGmBU75J
1AhFWMwWHkop5a1hQLpyyWN5Pvunvtwe+i92USjZzFD4iUG5SsQCb8ukJXhm3G5uLq640z3Bz8A1
zgQB29c/qpBSIjCl6gSM8PlZMd6mc7SeB8jVwm5pDpJS0K6xl/6/Exp9KBCR7SAuThqMciII5eQG
1BMT2GzCBP5sxLh5SX+KUoRuSOEJpUhwWjmK9cSfNNUm2Q/PBNZEZJ4jSjYkle0VKtuhbfMZqFGH
xCr0C0o0J2pgH+64jvJpr794pRF01DojjDkJptCK1aDoor5DqrrwxBjeQIbGon3gw2eggP+Y9kKa
IkYPauIudohThcFzrAoivfEyxwmZ/dv6Mw1TdmiMWHOpnWbZg8Y6GrnrGLFv7tqh3AUMs+Q0zms3
ew2l3b0/rYjWeQ9nQ3RYGm/3jIsHbY+w0RhTvC81YQvLtX7l2ttB5LClkeRgyRtEW1zaFN9XfCs0
f6MiIcKVlBQJP1AaCl1emn9/1t/4tPsZWx3/Yw8Ukc5wC8EHMIAf/U3gm1e8CcQAG4XjDdNEEtpC
s/Hjx3rW82nJBOTOVhdziBZx9EeCDor5jRJ8XJ7CCIgQNt7Ph/9GB9tGk2pwCWLxWRuBfyuXyA08
kOAnMmdIhhKGKjRD5BqjOuYcY4jTOM9dqIIDlvHLCeqQuIpkGxOEqxV703km8nPGPrpmEPt4tmFI
+Q6p8fBF9VjB1h+MS5o9k/06YvBzH8xT2ZudWNg8NUwPHV4MJyXxVmLEil1AncZRTaESSp6LYp+2
j+GDVhf2cb+enbmar6XpAPknn5RML6tHitfOKK2d2F3KdDFCt6DOXn+2zZC4qa5E+mbdzQywbdtV
9uLOnDbCHuegOKL3UrskAkIDUVU3zjheiMkkihY8IJom5v4i5NSXb8dKvUTzLqvSG9hVyYo9uQan
DBgf30sydJWkdxN7Uy11/2pZn1DNvfhF3RqJF9xLhoYQEsKMMR9Sx5Pc1BD+HlbNeW2J0uv3cox9
0kRlJ9pP/aLcacPV0eCFCvfg2KKzEQ5Z4yIJY9Fv1MxInQdG2Q9CLu09dXQcJJ0YywpafV+mYIzr
p4+bwsDwzsO8HzRHItamhgV7SKrPLFmm7JGk6rS+LUB4n1JKKHcTQ2GhHh5i3nAoEh0VCv8L8n26
jRfwsAtCpa5FzuWhumcRknopqF9NH80U1MEjzUt0O3Du/2ySFx63RGAp3i1ts8fVm/pZNos1y3jX
ykFvr/P9TgXwHSC0UbbKRwVs26SP7pLEr8AopyAm1tNmB5PrGVERcEsGIDJ0p1LD8Psk4WB7Zsxr
mBc1ead5v8DiLf++VE2524e85Hxepcmq5bczlBEQMRzyV6EDZC53jmYpppsJ6+lPAEdC/bpwGIhY
rlWYIBptAib6RCWG4gV/+AcPZXg8Kv825PvqRF6DGsL8TLwLX3gAHr4ZRwSiSRywScDVhTq/0roB
3tiVDjvu71MqDLNFo/5eI2GJm4da21RrVy03KVYa5RHYaXatyeiEgVzAJXjPRjDGrXG09SQInAc5
N6FYOB5Y+VAt/0RRTjucCmrdF1oSeht13Q7B0RamXX2fpkynEOHgFqcoTgY99X5BrDmemi8GlnuC
7e+++KajUrl6osqYhfPCgTxh7aZIwoapb6E/ZJgcJ4T7GXl38B1WZoR5WQrzv1CEv6bfPEMG5cHP
Fq5cHogz8kG6EPbjA29JNq+vBvWHwhngHP98fJIAg57PUccGVmlzGESA3vQNfL3XD43YMGVjuuha
63kvHHjAE7xN0Si4RQMCDwz2FL3BIjH2/2X7bS7PPf2W+c2AkvckQ9gervj3jdolaSzN0vcPPX8E
vtV5N89UZ4GOgFoOslyqCN832seOqvMKEnHOiPnEoLaSth8tJIIIwaQ+2GdStKiHXnFkqUmntVL3
iYPy0ywm90tKo5wd6TsQTyGfDhCaEay9CBT9lukkuDjV7MAIPOE/4mqGdn2n6TXHAjVRNDaXWyw6
JlIjdRSSHJz/KLr9cbazUfbV7fPPBPORDIvy7KH02ddhGAI1zKYbSlzqX5t2pBLN9zNM1H2AB0tt
JD4WJ1OMk9bPqGsRTXigl4Xqj0Lj3ayXzEf14ufpC/23IwGckW56SIqbTEv2DobWJfZDWRbmPT+l
0kt5svM1WHcGRanjjNsh3PETJrxzE67RBxx6CrL5ua7aQj1N8ZvAH9vq8dJBQepChDsPvqzXYPJm
aQ6bjXX2t6ceeNm5uV7Dr1VV2iV1YUTgUDMX4Y8p8W++VJ23Bj9Hkq5TFAlNKf274/DUZMIcvUMv
HRMh1vfOsYzoN1N8wC3QwTEIrtZwsdtgcYj9h6gp0piTYwWH4YXOx3N1jwduOg7wRyCqlgujM/mv
qpyInM34Z+9YwCavLwcF4YrJInw+JBNM/9xx0wSuQL00TVKPJf6ODt0p873b3x/s1P5551czUFwW
bSShlTSSMrGaXWUUxIGemUjLsv3Ykz0PI7WqBxSgj/N/yPczJ/fkDwLNim3uAxzfz5Lf7U6q0SHX
W6Yc1HtLUA6tC3dk2d7PwWQ/njDQ0wcqwPR5maPirZwUyTOUsAJlps4G0N2je3Q5k6hwtCohpp6C
uRpn0JoJtvN9cV05WurYteTb0TYtXm5nsVFcii2WbtzM7TEP/SceTmp9rTXZ6ZMQ6e6YDPFHqkZT
hi4DiG9SHC4EvDzlibWiyrj20UtKsnv7W3jAUcaewXLN2HZPyo85FfVO6UBiVTDJpOP0ZGsdlSIX
EPyuYU7UmWFij21K4dcWTrVnfw3EyJQIBMB1UThPuEV5U8yJt9I/JQZHntGkoja+QixYHVPNPiQS
iCLwfqyhwYrBHcMe4pwLBShEI3IWB9V04lxCZ7L89aB6I+6nb4EqdxIH5+Ly35O5qs9zXA9eNQ3W
xlmAE8YBE8506tZ77sTgQYl6NV35i7MqYf2JVEsqbmBMI8kcgvA3zDaBAgS4bm8NP63z4uEOS885
57VIuqrjjoySuJCUbyGqgzc2tvXahKqZQBQ31KKS6f/8lW9DT3k64fWbczNSc8QvhkaEFcrO6Wve
ToWs6+oMkPihUrV+yjhKegjii8jy5crN2ysX7WiAUIrwPjp9CRLLOtP7eTO/Tx5TjnF1rmww/xJb
gtHrQl3iFBRrOsa5q95FEYzWXmD2egNGhYcSR0kgg8OsNEJibcU2nx9GrHSpL/T9YL4jEpIcjrVW
NTAw6Dn/FU5I+0PArIUvYpSmdqMn56X7lCeREGfys5v0mJYxiBwuBffjZwu/YiO/1RfcjMsJB+U9
GZBKBaNRr6nmHNg/pIxEeGhiZbdDl7MC8CZrTJcutMLFD08wMIpTJWzE5zmz9tXIB64qcaxCYEH0
t30jaSYO0vJ9J7Ed/EIGoea1Je3dtCpqwoi3lWGii4I6zugDLN6CkWlMIWAW9hJEsIxjDTnffoqx
X0W+tI3IIG8vi25DGvhrs1hJZrEtxQtESGr0L/hIHh28gNzgiF1i52x79GBvA5ssTw2V8d5ZjB3X
I1QicZsIMM/ghI6vdCPnpHz9jb+kXnQ4nxwloaU29K7JIBNCaQm32xpTr/9gx1oe3gAu8PYp7XD7
bSRwurf3YeECTvtiUZ0v066C/zGYATEPhah4HDu5nxEVZw67ZTFkcW/8URK6ol03xbpveAZnjfGp
JiqDui2PZLZ1gGmnPjxzKV7nzFdSJhsYFgxIA+9eoAzSb2DkKpcf6JMJl+AwIN1Z/uhgN/D4+vnL
SE84/DKWVc5+gyPC/p1Jd0mkq6aaHpyu4Z+C2CxyGdk+g96cPAVpSZRfWncScc2HmSYp3uMK9d8h
zouWHcAliT77mSi7kyOlXiFK8pUGNvp1D0RT6QxRtnt7SIZ4NPYIE7k9mOVYEcinotCqWkuJl65z
hQ4v1c7/m3ll8l+CPaosh2Z27SedtmN46GOZs3yoEOmpOvhmtGwdivOfEqEu9egaQVtQNJBBpjId
9BCK1WFyjzO9QYQxhLP2sAeoNyjJkDs6jZwzihpRO3BP4IXoG3kKqIKim30epD4jYJ47VIaf1KGL
SoPDD5iFcw5xJmmQtNH0QQYFVXnXALCZc/sFspdid/12a0xj5RJvi4h6qDlq6u59qlWywpH9R4VT
IJpp4NbXg/FI9QC3N8vDnuATG3Ld55WkgzU4qNJ77glgQYCaUvxM4WQWok7C4Y71P4vgrcP3tih9
qZJlkIMZZ/HHw1DDikxjUXnmWuV9M6/ksU9xT9foL45uFf6jGluPY6a6BqnUA/weO6Cu5l7lPpZ7
JwTWynp+ds/v/hIE4sZTmwCgZctvoSAd9Z9Jx8kF4spZbWSUl2okk597LvCEdUQ0GBgI8w/lL/b1
U0YKztqqYMxxVKxcCl+SuyzcNxrG6gNWQyuZMr43ZCpOLpEvIZlBd6nopYEGgOkkj7Dg6VBWOJKP
5mjW76/IL8IuyagHSzI01SHBer59ipGjPSkFsDvJutvISos0N8jnvgD4rGfqT5ub8395ykvTt1wG
h74Jaffr0jYwubM6euw7j7eSc6fsdsXdvdzodtv9VZ+IDZn1W73zmqzR5iyTOnbJlbpHCUUXsPqN
cvYRHpyLHHJtOifWIT53wOrac2RE5chFea9vmkbDVhhMli+ioaRftaADi/+zfBLU/KEBEYMEJTBJ
22gp6/jvoiyiJPdoJULcY4WRfcaycHLklw4sZXSvah0PNo4zc6ZRIDslX9Uf5wyZLUh89EdRAUqU
dRBhOKY2+pdISzvouUTxV5yBw/1rbvru8iYoTc5HG2udDFDTLlBaCw/OmWj90RTDvJVhEpAFpSew
2YeB5ZacLGTsJJkOi0pj90Y8ZKJGxjXAKCfB/+0+befLupH6R1mS0fl0FSIy8LAUT4oYiJRiarpv
pGA5qo6ZJDG449MYdopMKkssNhw8+LlH+BecFazL4vtDR65diMDPDI/38ze2N/s0pr6m+uLs1biN
zgCTokbZYwmnGwMsW6z2UugQsJuXb+VO7k9OG/Ov6QfUm6APEmxVkU6OVceK6EKhM5lKHd4fdhS7
avqtdiaLX5peG7t+2g7rQAO4eStwIv+m3smjwBzNqzIN+o9GkvBOwLemYuZ45rPMknA62yP/p/oT
yXXoB5GpCt4GihkicyG5ZwaIstTDUv3vWm1p4PMWcXbCa05BnGX8xVJXQlPHGusMGEmovxLm8vlJ
Jrq0mvis3Whzsx2LrPfzd1KrQFHzxN3QT6Yk8Nw0r+ytmybgL0AQ+rOGJcQtQ6LnACu7V9NoPvrg
3EUGQ4f5janY4Aacv8s74FFGLsQJOqQEUtVqEfM4Yd0Ha4LAuPRBoIBlqqIUhohfRvbqFjQ+8wWw
Wjb98377xhJxXjXuasSO/u/3fp6eksdlMHokfUaEgez2Mdwzn7XmXDGI4FZzDqlawA2Zqkfd8PlX
xZv7fg6nDxdzykckNjDxOpEhPq7lnk9gDUjzkq9slcLs+DnFHQNg+mAyed51izSi7YQQKFSB7q38
v18DfQqGA8c5NOUaaFzCtrgujyTfEZrxN1b7rlYQYUmoz5LWWaJvi605OTGihqaYCB+K+HhJuXjL
gHABGZdjv1JOEmYpll/zP7FPGG3cTiNlK1SfgnPm6zqkRWDWD+CthKeQs4ofa6a6n6X6QDRbfGir
ax0Q5SyWahyKrPtjv90qUfwZSJlGlkISgvsiHyQ6NCSqLjm0P4v2AM+z+vnDLAYVkupSNz8yiOw0
A/NWymgibLbrWX1Qu3ZR+ufG9r9w+Hq/ctRS5KBM40d4FayAgfln5N93/V84UyMmRpBlN7eEkhDJ
sjK5c7WYuE3NWC8FAdEyy1CXtLduRYG6ntdvsikDu5rGfFOMhP4F8JX8P5+P59xgvvjKwwkHt7Xu
LpZ2M/vJSrqdj8rYJbVJy/3CYf7iFJVKxK3Q/KGogMDGeZojhcRHZNBqLHwwsXkRToAChIBKmBbv
44+3gbwd/VsIZbJDG5fQg5C11SSDacxveHUZv3f9/IpxysP4jUCXjgXsp3+nSeOvJE3cu7eDnm6r
jfFHhaHuy6HG5udmByiZ9Nk1rdHKHHxogf5Lj1piibL4PaRmNnwOECRpjez03rNHVdvmZttoEpCB
NV1beRf5tEjOAFyu90oeLRlmkd4XmqF91us70/JhcALs0kiUkxD07cbqkkMweofEWigjvD9dRpTG
5n9DDQq/QELm6vbdG1Uj4vUcwJ5gPwDuq9N1RLEbHTsdGf6CKsuqUISXKlXgISidrqYdbH/sDkHn
bZEtk81J7L7yqmmIIn99V34VhBruSZIGKd9tlIs+zcKhrlGzC7aqGpI82BF6aoNI8khTN0IDoVL3
4dB8rE9VK0zY+6UiZ+/3tv9mZjIVL9uQ2KZwpogMlCKkw1e5C4pjGMHwxTPT0tfd9jYIRII2S02P
8p94EUOc1vwq21g1C7h+6fXu8uOOj/O1kVrqFTir2ej4NF9aVdXvImJaEMsB42OeCkSOB6+qzHaU
okkXEJflKday+4ojxAvdwxogxvpiM0mSevESPqhIna/HLw8D8G3EKl0xnCVBs/U+2RiNLl1heyy2
v9BICvKu8/WeqBzk3Dek22jYVx9qULMK1FnBfpnhhtHh71zcIiPRlNCPz97qn/60unIf0qeopzJ1
SLkCI8SrDJ4NCzhEdVaYLfPKNpxonN5UHhehFhk6LlDEO8PXIrS9h20MUkrJMcB1ucFeGgiMq/eK
HY8gebPzoEuABSRLmwiCSbXzuq3LK6me2tE35h5xtfTmoYI3TMJVg+4rp7DH/l+7xRMgxQlf/ChY
lK++4PMG1NvRYoR0yhmufLs47ZtQwuCwYhgOnQX8eQ6mpIWFiU62QkQcNs0yujXZWkrh+Sc/BXnK
713YIBmnDMTzdrsVuYvrzug1MSxEt81NWVvnIdYghZTUmt1LRi7kFa4z06s6vuSEDRWStFkICc5F
jAUsGpnf75fOGMU6FVaGaB56nWCk2m1RaK73pcZTBC872dnyermwkAKKy4G4EquN9S6fPzHXvF0s
UMu7psBDBAF+GU/bJojRQEiwtMPJ7J5HiQSzPodOyWSVFUovIXYslyP9vdZH1bXVpE2vyVBk63kN
XZccCxcG5mrYKdlOtGeZ0shxknUMrNK2IMRtLNyGP4lLg3w4jP7xY9ytoJvTEihXoBKLd1e8Hmr9
lNDCQJWsFpK7TZSEKbWCPFoO9mZo/lvLqOJ0ZSd3vLkmdUNFe0+zkeqirPSPl2/fMuJmwcFESI+w
rXzAyENEu3ePHCNCbjEMPBRjGD2qC9yjxn+ues8uo9gC61qrZw1KT0mFmyy79FQ7zh/0DN4eRrv6
udxSSFU6JbwIlGnAnrIqsYYKCbRTQWbDunEhCkFq0filZ6tl7adFCdcP/bTcG+N36DVaGnMaoh3N
2dGwaGxZRim3Vul9vl5V16D8Wnr85y6SW05AKQSMDTlIGft1F9S/ViLvlm9NdgqrZpfvSRysSRJD
l8Jpgp86Z0S7QYrgKy25UiKZzNn+wYg6AQA0TrpanabOTKKJ/smL3oSDHynYp1GW3WveJ02kqqLQ
BejkEK6T4rskO5N4E6rDooHCQInsVsbLlnQFtS5uYb1nu7RG9H9S/gDveFuQfDugBe2PzlKpmQje
0cf8kQI1DkgX9NY61towUH/seChkGhcjDjyBIIggOY0f2sxX/1NpKYIGosGGVIXBHGwdWd6v92qc
qkBJ/+Xs9XOwXTIHgzNQHgni+IuKpcKF1Y4neN0nwiy7ks+eqYc0ypykkVU645yJh5T3fY54O6C6
UXaE5/AyTOLtD4y3Iwd5IMk+oE1B9TPxIJ7OUE/dJGupptSK2Y+3u0u6O0qu5RAhy3nVvEgh51BX
UjPBomvrkdL71tsxqwB2geDN+6/XnYLuwtTisO0EBYIUfZNVlx5PWO8a/mV8P5jpzyIWWyEr/oNL
ZA0WQsOtgw++b+pqbppvIcviV4pzQ8ZqGFQXiNFo/wbJsFeTDMeE0chGDrTaPnaMftbKHxKusdVC
6nkVd0k6uukfJz6ZFMWzbtquB8QgqaAWPsTnZY3o5rgofjebw9pKGWSBToWfsIHeHKl17T7nIIa0
Hsi5FOoOCFctSsGmpe02KV7oIMiyI7f5/ptkoYxHS4R2gHD4xp8Rc1pcI16AJnCCoOBr7NuXdcKU
R888xEQ+AzL3AzPN+GT8xREb60lsUC8NYnDkaGySLqhlbWXt3s4fXThhh+uU7W2QEz7PMNMAaBkO
TC3lNsJcOcXvkP/eBylWQb+5paFYaQtjOCUjAwfR8KrFgrqiBCDTa6CT+ks9Fh0sIBNwej7xd82u
c8iWU1Im5DDZkTLutUBB5MBzS0evPWPN90YK9lpJbCJdM6A+KhUaTaqzShcNe5bVSKWMgIP3Ufb/
0v7tE9TQhSG0y6ENPWiRaN5G3s2vO4hmg8k+0oN6YuAkO/pJYfrdk4HCE/WVpG5oB/pbfSBhJ4Hr
koy1ntppVUTRCTQsWFGUM/Kvlp4vAq+mPE/unh/9yp2uArMSmdnLav+7BgtD1rmjucRMOE3kFIqi
WceFjKayUZX8H4t2+hUhBT9AlTAIIshMDCBCLFbpy5HYNd2V1oftTFCc/nkyUSKSa4eYVv+Agml8
eILJNRVVtIBjMtjuBqSvLWffmBE5GgGu+jKanng+kFpkx8mMfzotcVXposE8Trgk2zxQfhk1ys8H
7i7ga6ji9IP9jVnivAenctC+wsv2/cStaCA9CedifXridoQwj8/9Cng8z400UaN4BV2i54DWLs2s
7CtKAidYlgtgZptbdBuHqf77lElwWSJxy8xO6iNL7VvM9eVT0AXZTn6s3920CyWeetRwYq5Z9Cfv
6jDrnpYdk1MQSZjzOpq7CIKepqZh5XjqZaqhTAp4Z+NY6tpqnzXNMYiiWyK4hqvZsXe0L2vHdJz3
KYFbpBlQV2HAsLCh7l1jEgJGdkgFs1KDBRmubb9VAA+rONCbK4p/7UZzBO3n1hUq+YzC+69QiVMi
hRBA+VAYiAw0HO6aMaL1YKPCQBnvXEkvLWZKQWuozn/yuAoRkieQLYErVbQK3St/Ov9Me8wdXP2d
GoGihVVpnaiGanNHsHbZzeNPM1EKZmPguQS9eRZ5816pzgzNwWmMBZtXQrTaPtA2zxy3vZ4/ot+L
cQcJ41jSyJJiWtotwZbivJj2vDjNJtOeBYIViNMeD6GbhBB9ubOIn5NtONRcB9L1icWswzBGTh6J
ez+S3pl4eOzL6h7b3ryWpVtYGx9nZnZytKQzQmQHStunluuCk3hJpSINr5/Pfvp/cYJfzpIMi824
VoOUWD0FOrBswAMim5MmzrJ8Y2JzwKBD6tmB25Jcahj378IuSkE0LBmS02kEhXVmBXMAD6WuXB/o
d7Hr7qNH1Nn6Wr01C3khRepy4yHUFGFbGhxwYsxwesRx/eAqPlG/RGN8FJyiBxaB9ggxHpqpYJJq
AkN5DO0VaRpCqRYbc+TRM/W4B+4C1RgrVOAYyaXFMETtHdt6hvjjrxEtqYwSf424kvlfwT3WHr3n
4FnIhJHnmuuILZCCus1yUdYqyl52l92CWiOf38mNQw2iEXG/6relzow6+XSmwTrHCOdnt0Rt2FN4
qf8FBfog5Tl6tgKJFL/Mj9M3HZd6IlU/qEkqUtjFYF27n/RGZXxzE1xyPFRqOc2+3FN4nYPLE/v9
6KJyXB74aZNnLCys/4f6qHL9icULl2erixUROS1oVKf+s8OMPRiuIITA1/Q5HIxXBDmK32nv/IZV
N3NwIQqiy0XGlO9WYoPGVGNGa9nxZd4oNBzMI3njSU8vhfBop7YFoUE6f01A10w4jERXykxvJY6k
nededw2RRWb9WrOdkh4cMlvpDNoDPI0e/dkfoxl5nJVvsFX2NsnvM8UijpAfjhu2rl8mBzVPkjaO
14qbQ0DCSlZSI7Xq1rKHZksTAvo8omZawEI6Lb6tQhlrsQPsDhVQSvfKtvmgMLuMpxPA9daqy/5X
KGIozIwb9E3LfybB+8q8WD3Qr23Bzqv3f7ie1cuq6EPXpRBIh9Od348RJi5adZeu8Oj3tellWcqU
FzOLB/pYRbg0h1WL5SpxlIBN6L8A8j/veRG4ZO29NaYbxT3Sr0qIxoanA1JbqdOxOkm9rQIuBefn
aQQ2Lo5BGFT1Qe3+lHGsG1sftHdNSjolTEREFQDna8kcqRCwTLe+oD0rrIyWsBFVk3Rdimhmb0Fz
oH7HToaVr+HAfozD+oiqz4xkOEa1qf6TL8yl95X2VaVsN/BLYWhsUDkbCJXL0JlKcTi4o02kbXiS
v4VbOp9Do4SX9bcY0QxWGKde6J5Cflm7Hihdmw94k17XM9I/1Zst5wllCwioDIbCF6mNg39XRSqv
fENOoGHHgH41ASTl5DaOpnku8cL+31aq7sJYemzpp8MkunDNpOwa1jAGObGlEqSSF7qVphZp9PXk
gRiyiWpX//nTrk7ce+qbn0wMhjJ3gps76RGEClkHhTxX/Atrk7AUragXq2qUrDa4LqrMo8ZHv3D9
88S8jRoOZWkyKVKrgaENGb+COCVRIKNC8LzDD1G26qHSSbKn0KuJFe89rol56oRGfcrznGKKd0y8
v5+v96bKT2ip9QEvB4tUrsvgiUaBF49H2p+FqZmjPxMepbqedFRxVY3LQLwX5PRIuuzK80OtTkwo
JjwZLzrYo26nEl6aZwIB3SBgIgGe0DFS0wH3FpogBVaf1TcgxkvPoRrAFyZxhkk8zjBRkbNcIZZK
62F8cAjvWdMn56NU2MWP6n3EKlI/vj3HJ92bM+0xY2DpeJDWESyZfrJEoKA/iP9cONaNRO/UOCOD
l5w6byXoV5J9eVGv9WemFosyZoB3AIvA3ROYB9m0d9tvdRDc8sTETl3O821MPX5nMp5wOyzCXNwI
NyLDUq9Si81ioR8v2gu0nyUYrZvONoz6TzLdFrI/NCTiJmaC1vVWSjOTkerqcKR69/AKtkj43jBU
bKPwWPVDn/iqqWzfK79I7BTVc7kMEnyxc+fOt92rUuBP58QHjcNhx7/mYadEEvsCGD59Rr2DRUrk
66w0YE7lw/QSq5BaAHQQjKY0HrU5pKb/6T/LYivDOxVeKnZkrE7lHLt8lX3AxxqErmVSP46mSprs
ZvOzWSz0UoxaiEUI8qrNKNEchY48lxLwfEVZV41kQehDcb58cqHeM48qS3Hl3aI9/b8t9pwZME7R
st5kBrMt5b3iHwIJ3VINi/HyN6xDgr2ltLPFKpHBlt/BFb+Cm6rohGaqekRCZns+U67TCgXRUuhP
zs0jWZ2gCLMs6RKLXhYpIJk0VJXCiikp/KcwYzqpYyo5bXYJupEg0NywFbVJcT9OBwefyNOCjRJ0
6dnFGNs2Xz+pJyxWFfC3J59kl2CvigN/MUeTvQoiSh5BdeEO9j34SSzJqq0sl8Dxa9mrpMs8n8Nw
geLh9o2P+fjB4QGkBVYZI9YldJyTkEIrcnK1WHZnPtX8OGrAFG99AMQkVp5ZRl3jq3ftFDArweiI
VpyFBCAp5KfC+g/F++K1PzPo4OM2vOLbG5Ce32MjEJ761LK3RTq2tXThCyZhPT2C9DxvvrqluSgJ
9poHNlg2DzU6+bgLx0NmYDNv9yfsFZgqcp9gPO0vJ8zIVXBlcfft39lQehrxE7IMqmi9FaH4IDrn
qoxPQW+BDk4477EusKP4RJlgGGtRSSwSlo0k8SdhxwKX+qPDuUO9glajGD8tVwoJ1miJLPbZ10F9
IKGYkIw19ypege2qkTqYCzBiFvsnv8RxmpjRq/xZBeO69HX2Q5l4Nn7KG+tWbaW3f8cbAvHJFarR
sweev34+adczKwt9WpSj9oELftvdQjR3lQclN4gAol9LY+Yd5fwf6wzeiq5S8OPPwKdDQtj0ff9D
edgj489fjcc+ZZ2Rs6yopX+Rd+WDGaVxhf10huPKgu7ZjDOAx1IlGRKHnxi+n+FRHIN9EHKEqAR+
yVis4wZQdadojxdjXUvPddhRsqEyDb4mnFcbHiip2yHlc7eTB3M4SDBxzqvknlppkFvACumGy8TE
LW39Aztkyip+i7L7YA3guGI6Wc+hRpuKL+6gYOrYlS29wCX6pzeYWp35WMxK4vI+mwnROoNjYMZt
Ywo9PD60Sw4W3iTEpZtJOdT5HUFm4coHHKWcUZO2VAx9xWyEqKnBEDp1U8Qj5H3PacQkijGW07oT
vih/v4+xK6CNRv10ES4DOYU5iGD3zMGz2aAjRCVdVGNJGpVpmrVTtAP+Bgc15dEtUZE/20aLzl/o
JsGzypZxK2JiHO02iSRmy0DPVejnazVLi7gq/8WRLC9A0m8yvkXz08uUdrHw0fVLqKPh9NQhxPv9
1htqGLXDatLqLl7p6oMR//AUe3QC9RQGYZdJddOHKxiFogJeGF3qqJ7TT83Bda0EQOPfSwkU70fm
Q3LURtvgVlg0gU/5llS9wlVZq/kAJIEA0J3/0DU6HpkIJ14oEx6snQl293fjCQgS4YG6YtcmZgXZ
OKgY7sq9+JQCu6eSmeZXYxL9MIdXevmtLAFVCkZfuMLDjJgXgm2QEqS8i1ez0CCmLjSvLKwrSmR2
q2/zOQGTcNOW4d0gEtvzQK5chhTruZqWcbGxkknsDFZrObNFXSaAMYT8/hAJJJHB/9vSZbA/x6H+
ONJRfkKlb9Ph48arR1mh5MY1Qw4bagMs1VwIgTvefi0WV1N/9iPRxcbtQXCOofjeKIYG01lVDP9C
NKfAaarKLNAcdtys6wcNRmNY736xrNrwCwxXiHOjwQz7MaO278tB84FK8tGFWVpwNd2QOiiUwFto
Zo+Oae2T6kBycDFyLgtlA1Q48Uw7AE/E6Jf51lLOz2c6EuXOAFTadLxcRQSKFmoERT4K9etQ0yZZ
FNUVzHdZjxxr1epYexH8M236BEXYalfaN9vtFsT8vGSqzrq0YRcgMP8M+3eXvZlpQ/+czJpTuMRk
i9zTbire+MfV1iA/pCRcP8VwK+IodRE86tV5jMftEOLegxdC1cN29U8tLJ0q4I+xAmTWAJoW3rfU
zabt3fH/B10+AMsTU7lgX+qkRCGqx1X33P23f0AK3NutX50Cms+UHrCvgY2DVRx2Gmpnr00qjErb
ZVEvxqvmbehiHgiu0zFDW4GgJrtiIWRllEF8nAAjJIRpybvsD23+4Xe7uKe1ThbS/Z4htOunKtwH
53KniC15T0XlK2mpIm1MKhxy7Xf6xV+McvC9hBAUmvQtxbli3uJkReXjSmFzmtNm6IGz3/OlStUK
yIAd9zKw3wpCBAV0e/kbJQoY0EawCVByIQKsyL/i2jMVjf+IUOQ/uCMKH1XWu4uxYYw5ojXdEqt6
kUxbcXxYXWSVvwtnfciqCC2DioJFOM8tLaN9CFCWWMFEIpfFrN5IEGTR6J5nTfKOt5WCHOpTC1cC
HYZjUHWl0JpcybRa3EEqWA2hpZakxr5JxAWvqWvwmnKTqShGze40SGWZYfLgUPp7b6k0mLzwMbY6
uv2BzzgsI+gXpEi6sgQc+T7wF/HDiVEBx/N8da5QQzKNOb2ktdGNPEpTyXAjXzlOF/KL376lXS9D
e9k2yWMOmvEnudA42JVGPRTNVMDtYjbUkYWwkpKb5LV1JsWtTwAkYrtJUehpoEO65y+ohErP77FG
O4g6g1X5994KW4VwPjkUGiRBK9jvmuYsipvehcKDyhg4i6ucqqDGsf9OlmIYKTL2kYzDiRAVXXpP
HAjhR5gMdM0QKUyUCYBJVs35FniC/3By9al//ZvMTVt35NlLZjkPBubeGDGvp4I+DIQ63wzpAvO2
qBh+goEX20X8InJpIsuaRaVYNhKqSodKzRW/iyIQMffJK3TIDCP8pk+4bg1swy9z/n+cjwFT1Ml6
8equOIslV0/56t1wwozvc7qvSD4ygUMUD3Fp2zr8U6RUvLMPfsbDLF8PSNEQRulqxGdB6Sq0fjZE
e3HZ9i2llPcLsQMUW2QUZR8HS7NGG5Q9p+JQgylYE0i0GEkwZNYP+c58ynjXZEVh177I7Kc3zj3b
EbSbPKOj1aDBpG5F+90v7+d2KajeWcO/tcT29CTS8NwGsDBXi83mBvLqs036hH7VYzHH0xDoZPSF
ihQNRNOUTJgQTxLjqCKoRCF2aSOFC+2b+ZaxVknDZA+wNv+WJej1t5ht6nkls7UMM93noIc/0DiI
j445oZS3TWh8aFiIu9cJ6SGbT4OxISo4pEFloHgFiJjViqtLFRxOC0t7mDw/rkrNwGPNZjBJP5gw
ATGS/fe0vOQy/4tkYba9E+Iv9iYHHfaw7L5df66wXp2PtEf4VwrTCRmL5xmP/D02R0aeKFcz10hK
ocR4uL2UM/5D+9+HmmIlaIDH5HF9IpxTdRw5kt2Q6Ah/y6e9HQs9dFYn6vUpGn30eo8vAoTwLEcw
GCQfY7dXqK0uIXtBERTlAPOvrOePDr6LHzI12kWEFUyRYVzvJQWCK4s1d2+ZDkz0lVlQlN4dpC43
QcmtVXOv5clJ2h95R96+yZB9JJdqZgPvHJF+0va9AorLVOrCZTIlV8gUWv0j3KXR4wYbgb0L8Ths
Xi9skHp8t+u3P51FRtOSFLAgIvmjPgKwoeOjNNmTzR1t8MLPRLPOLiSZxQNb99MU/rfmthJdfKgJ
/QWq+UF02JHgJki128GzvPR6hxYOT5Bth/GrzG6g6BLvjXX1z29EE9WmbyF/jisVmSffBgPhSnqK
ONLSARU6SApdOspUc7dkUFEPo0BwJqSaZj6E7wvDx5MU2xUjVKOHD9SeLsXIbXAfjWfs7Pj0pU2w
oJeZJEsdERWhCbLZCZHsVMkC8PzJo9+06k7y67ORZwnIk4wiIp1pyR+JJpP3EjjZBWVOCZwndeRm
i2NdJlATe8dPp3/8UQV+6eTXUokbtL6R48GJN4DQIO8zcO4gpxLV+hurSTphmMJb/iy8BurAW3/1
3taVqL5Tw7+3xyLy8EOTT8uprfBPWwzBEaJq4//A4Om7irsbBUmUQ82CNQMigqFFZiLDIkqtG9Pc
NKgd7ziNThHMR84oFWeqGFTmfVhUUjPBKoq+P7wtrKRw30jiHzqt9fMtegn1jKqV9/3fv5WCTGNF
YtDYwJX9TOyFOZwsXMl9SY5/0Gle4xqJWyPJfPt4zqBR+RHkcghcfZdkydbO418p8YolehmOaUM8
sXJTn/JzbFpmxmBBGvMNTUsXHnIczquqA+5U1jwUGm+tWejbRXI9GVooJkUrgO/na6c8RTzNJ7ge
W3S+cYsw6YFEQ7gWdVb7Tu+8tgrLEYDYn5fo1mJYMCNBqgw2d78yeAcYezRYDf+F0f8A7Sa8sq4C
Y8XeF0lidxeTKbia6nTl8juviWfgFjElsE+69JXXXypbJ/P78Z8geYjRKC+b49zUjUdnZLGZwyTW
UxGZ973/4SaFk8yIRNxtlx3azf/viqP5SyD2CVPZAtyPQYlcvu8kRrccgJh11jDiTIUiHJ2N2dgS
2Lu/o6XRF2X9Dn8kzkkwhRMaiocB/i94okWHVfSvPv5Hw3vxNXfuxe0o5A/FY8SefHJyT+c+dh3H
BcZbSHfnGrdBcJXSYGWFwVTqjWm3lbKmZULV/ubqZK7/w2kOkb5zPZbMq6JHN3o9spwV+hEzdw14
Qq34NHivoN0iGS7USbHMLG3/6qvpwQIdpDwjTh9EvcTlhNNN2CtiYrriCJSVQt/SFLWDQLbHAF/c
azhsAr/hxxXWlgzTE6ktxzXwFSR5iwwzyKoVjTUSB28xZ7J/XnhOxrUfTwkJo9Yqgu8p0FKJHSMn
xq6ivwA7ZAWPZOW3+arAxtKoBw/E6O3GhegY0sHfpwJOVnaqWmp5YZzo25HfIsVPRC/Kbc8zvxyp
6RBO98Z17EpkrHb4W+F4osayYL1lAX4pi946lDvsQzQbWtuU48eEeZp1emLH9n106Eezz2Rqp2IV
uU+J6U5qisbEdVf9hLIFY5+63SHb/npuZERH7MrWcoxgq6MhjmE9kGDjYbAcrJIQQQGkTSQaHFdR
QtVd94go5JK9Tm9e/1TnUHqn0FypF75vmsdU9rAjyNHYhDF9HMAiTCCqzyPDxOYY9AQMnjPmYXfs
7b0BsPmQw3MkoJwrq+Te2PpwqUJVmSpv/p3Z6xEzakdqsMimQ5End8b0hbY9nzBBFM14d3JtOfBG
Ye186n3ZK9A8KvxvX/aOmRZ6xrgDAHwVbIO9oMGqCyJ5oF1ccnXvm4CvLxm1XKNE827lHO23JHOx
Oqy3IxPmw25NccsILdKmNuxsnL3S6zM/xLlq3IYay/hfyWBGlxslCgvnixUj4pmPeyTVM05MT1xS
XP6NJw4yyWo6nwBcW9IKWBCQKljcGs6ZIkYrluAHROMCGOW7MD0t9lsD5or3S6/wRE4PPX2GQUzf
o5QINl/FQs096Pd5KIaRVoxePeQH5u8QPDr6v2DKJ6VZmIQ6YJx9CS7QQYwM7BNjFr4LC7sAfvu4
HEPj0mE3d9lNoAaCFeaj9DyfNS/UaZ0fVhHLqFSsmFO6F5/oC32AL4HpTREyf6rkZ5yzzhUgKt/Z
vbsj58/Bg0VD92J3rE4J2h2aP+4TXKibsb3DtOAU1HHAuQuNdkujRNx1P22nPU/O8vj/l1y21WzE
kfNEMyFzHWLTiWaKZTaSQpkzUXynv3bgII14tRu3IAhLTSjkicvEf/esWoMLzN27JLvqjmKjGvAV
DMrVK/z7/Q+RE2Bc6cKqJxQ9QnejnxeKEBd7zY/RVs/BOpFzxd8g17bfQiOBRVTj5xlYwMd5sMAR
9oBhXA3NbtHrUx3mf6RsS7gYDexMIBJpFKnXiGZMacbgO54p9OLjFf6yhRrfMBaggNUuhBCNouql
O/pyqZqPsifJAu+Usdll3J0n3C/YveGsbOl0qaC6kOPey0N0SLuOXfUwq4BjukdkwzSP/OZX97Io
vmtKpN1F45/zfh9ylNVFvRNpCqfD3F6ORz2bXk44VWp1u8puCypWP8r787nIyYq/La8O4rtEHLz5
h4w81cMzJxzhr4wHmOVlqngXZb2wggahZtZSzjSAPQmlqJi0ImCrSBUKfiQugVT4vhq1XkDtuNO9
lCfxpck97Uu0i6QNH9KPoKtbz/qKC1R72dPK7UViFGItVlxdCqPA7gNc5pZDaApKHTF6A4kfwuNc
6LTHA5s07KwOiOZLEc+44Lvl7wte0n6D9E9f4tHdrhd5yieykKcRMC/jGgicHRII1UhgKiKwGKr3
CvIyFSdlXRBg6i7TCQZYrWvz9zWvmI01JXGfovw6t3xK0VjS1KRNwjGS1fYH5dHAe4ioFpdlHD8a
ZNnOim3PnMXoxvRSvUqj+2iFARfQ6xKPlKksAl9fzocmx9145eAooRaGkY6EDMOVn+yP/v7bl4ng
L2+2PH9916OU24TYGttCAdaDifhC3Y59vwHdOdWKPXPpXk3F0wRtJric8heGdVAZyhKvibLkihDz
gYV5yO355ECHCEFwukM1PNiSsdL2CLKGPKoIsJ9gOk0BtgqeI4AOt4bHlKT3AD6kzfEMPY3eWXRO
M51TMTJUkiPcH8Yijg9tX80LbKaSTTvAYTGgnhj2RO/kcK3QAOS6981RB/uYR9MK5F75daHgrA1i
svpaWsE7WRoJ4X3gk+gfhKenwXeovNkWw222JNzVGdjGvh4fwa/ZLLGqiVv1Aj+W/62NIvEGIu8n
5oBlaOovwlDOAVKhP79/ImB3f3mmFJodeY158nUa13Guw0HD8X4RWAlkd9npqSN1sTRgz3cUSK1z
O8L9g3BZSi9bQUGoAjy7nQ/Pzji115klOPH1sevlW2z2WIxPDGqYwq3LJFLRPCoSG14bnQqkR13y
c2Mc4VA6yIhWf+265AH+0+31cVYsxGbVhAp+8Qu4nn/8NUsLnbfJWGewwQJnuTo6AUiIm1u9vXM1
OYAF5DjIv/UML1zFWNw8Tb+KYsSy235IZHrVKCHeAXnsmce0OV/a+thEHKDUYbOjHYx/WMngpMGR
sEtyiLt8NOXs1SWq+fd4m7QsCjaxmnKQc0cIMWbBYxg0PCoWHKz8Ogt0cJB3PdfS9KkU02MevdOG
gxU5wsrnh50pLul97UcemFEF0yVozG8qo3rOTrwWTRwEA8BWMMSumnSPUS06zWzqgiUqSIM4s1Wr
ejNhGXYgKBODO+4ZsOPfGiSeMcf6kBfqCS3SFbBBwuoaj0lo6AUOiQ8F69t7ick6CKgwMcSaGg+A
mH1ZdEdO0eeatp0MWz53+2Y4yvJZOfe4FnD/l5brOP5ol16Lrip02S7clGi/kdiWeQv4fWaoCvE4
2asoOhIgARzscGGvz97LoAaezmm4/eOUz3V+Gc+RUNPCS1rDWVyxv1MZSv6tyQNowH71frjUCtK9
Us8dEHCLfMnTPpBCkKoHwFHCuG25LC+SlE5BVc0QN5aR792eBlw/awq30GCc2YOYtAe+FizT47f4
/7C9fD0UCnKSHSY6bCtzIKW2g8OtlDVPZQ845l9Hdfnxrsafn48G2eDuopiKz020d6vJfXFBlQIG
6G+T4J5ZISFkRJxBQlWjWNBfenGQt6BhkCBKDm93yojYrG9aeI/qvorbDKMVtvBFTmGNp57Td20q
AOVYRe6NgOX/UaQBN2A4fOOoDKAbYK38IOWnPe/q9mynaFiDN4v/pF6ikwOlhU2bwSosYHSNGixg
Rd6+1wf5GWVWmiDwjeesoTGjKCh73E3OSYu8NgSskQG2qaR4kLlVSpNllOP0DBPltUXuzE9lRYqN
ucLjx/kLCgqH5XYaxF7RmTjntaMCZHUAt1dIRQpTrDbwhxGBQS91TN5rIARAyIa5f/Cz3k+8qEQh
9MxsDVIqXX5dmhmHte7TLaN8c51hWliSYm8vB9kbiOAbeZCcmfd5hIjiNU03/Ywx53oqWWCoixb3
OxDLWATpQ0VoDz7I0+/y9zELjVrvsycUZPsR9XXem586bm6yBgNFzItTJcJUXG6yrOsIaBAMJykE
Yf2uHUEa/pPO2TKDldCW5M67HBOBzsEvBCSmAtz6ifOUluxnSlm7avlEnZffFp4qA6od5rEfdh+i
mvtF9FtyH0JsEdZWSuCIyaVpmtsQ7VZI5JcEs4+/ZTq3uhgzFyC76C4Y7dMvvcHBX3I67I6W9JEW
KSffyIZ6Ll5lL3/fAmq0PWjw63opdDHxF1q1txLwDuA0etpvWVYtiEobN/PmHFDZue3e1TTuKa3j
RMLUXnrXwAnqtiXCJ6h/v+3dWlHSnxH5Bt7q6m1KZW/JBtZX2hgLN1uuwD6j7HAk/YDi04Vkv0/p
Sw6bKwo5UNT8Oc6MDMr+N5F+W8DihFq7mGQaBmdL9C5b9oXUjmJ+Tty9vfxgPQOMDh/MpTtrSRnX
SFuk/4b4N+vGE/zD+tLS7xdbSC4+OsMbeXIYGNyGF2wNuVjjHVPCeluh9VE7Nq2u1bUBNaKwAR6K
S6/ek7RRbW++dLJqS3IMOZC9KsOTiMmVzOvxxMEWhjockzNg6IvTBouBGbWPxNboe+q98Y/aqBJV
235UmVX0MvNR+7cP4BooT8xosNdsof7ppiP9ahl9VyBhUUtIKX1XUc+ZdYrOiBd2RGpdlp6t5DUX
UtgkSZIm7dq0EOl4XkZXbEVyC8ycuTJNby/FdunumSv7Gj3UHkq/JBfGtf9Lv9H70rEsf80GD4+D
3WbyrRHKzUVNsx942zcCFnjh6HPzGcxbmBboIZwshL7BfQ2zyzgwiw3LyM9v5p8YNVvSrqzYzTFz
Tx00DygZy7SZQScu6sbsoHigz0PU6L2JAm/+Df5tBH1eKd0D2PGz8G9rMmyQj+DDY0VslXPCNdN1
jfeXH+1QAHkhIbRLkpzp1xeeg5t2rrLkpeevsx1JqmbI74gbVK7tYLzC0KkRBzJxu1olSz9yPk3d
n85xo1Lm2rPBbm4cLQn2O640iiKNMbwjVV9ykrRfHhB8dd8eWXe3EncDZ1qA8ioxh7YD0BcCrFuN
BkGsNxDheYNPhTe7bSYF8u25YgkQrL1cnw+yKiUVOdPKYp8Rk6adCerlzZZWz8A1XJMBW9W1kn7W
t/Lo/166fZRm+fpMjZL6HaN3JMO+mb+bMBwBi38xALWxW5CJHhgKSSxcfoCUfpn64Thky3GQdvrg
ZBHXyoIT1f6KYYvIM9wElsj6JD2bwPfcnN76b1SAyqYvFxzd/7B+ssHJhbTAQkaKy+mx+PWzmkTZ
8Ftzbn4PNSaqlPShUQf0JYTvMnEEqldadv5zoi87LCJS2dlfcbxiEA1LsK6ilI6VdyAngfg4gj2T
+0OPiLe+XTcHjRReT2eWeCTaphzkZBSHSqMBh7v99cPiOg60GtWBK5qFnE+NwcZ98G1vhAoV8ob3
Uk9Fg0CSK5ahdmZXvapK7kR7sN0UYGXj4PXy68r6mppNK18+qDF/wpyvCyB6WMn7/C77A157VRGv
g/gYcIeFtegOwBIGKbXoa8msdy7ermWZVgSj/f6ptuONpD9/yEyqmDTTKpodVAEgtAtzWKh897Wf
PbfRZzg7akI29OwcnnDnuc89LVNw26pbFZDDsIFq+S3dhKL3dFL7d+2U2BeKYr9MnRFEMgCjj+lA
MA4qwx/d4x92CTArEJWJtQpDPoE1GezbQfSeiGsnOkvL7DbQ9qT1V88UXbCKRRxFM6Rb4DxmtiQT
Nqd5HTBTa6rNRyFh1cS6CVwYflIKYebkKqbMHZhJghgF0Hr8Tc7OqeSfCKRqiB3+oTo1BuJDDLrI
+QkTzZKAg3M4Qq1q35OhwoRDGDV7B/78dixYdXoMYQqJjgRu84LrUKTNkgOE4ZRkAMBWUJvwyJx4
lIL16hnzhM5qlB+CzRnEqoVsfHb9eAURpspn3sw7tJVR49ZGf8OCyiOKRrJO0zWaswCFjGQwIS4b
m1CuJqPCzPEvXTyg3PcLx/AWKm8YGi3nevCzyi7pcuNhyrz9UAhqoNHmdd9Zu2/Eg+XVY3k+Yabt
UrY9nAuRfvQ2ka1w8SVaqFTUAaLYBCTpU27ElvVT8zSuCsZftubhMwlT0G2c+p0X8ZqPOu5d6fGt
Zb5xuPwa5MeB1vl2BTBGYaUHp8OxlRauN1LQ1fKnNf5hXK0pfhxPKBqdwxE1Z5YqRU7fd/Y4k5Vg
NkZGMuGEPHOl2/hopAYJGuVzuXyuRo6DtmyYY0MUFBkq1cQGyR4on29DnNDFs0/OBC+8FDC9OaoF
JsGArQEk+raCEPbnSlNd75FyZjWABS/nDW0UZAJIFv0TzNP1zzv9juTkfa9mqVIAx9eBcvKMAg4k
kZ7JLsJ8JHAkY+QMqkTw9H+kUkZdqcWoFH6tVoBJDmreFecsmmafSziv/YgInrNZXl6x5nVka0f+
O2SHJBgeMWlDeZRCr8KJocXCrsq8yK64DrTBxtXe7pcYOBjGs+WsKNTL7Onml4lyD/eHukjEWu5z
XRgMnHuth7KtEactKcsuCkZXIY1FNUVp/XIZYJ9auLbuzVPWfWx3wYJrxr+QUYCD6QbTcKSjDPrr
X918obM9kVCbEo9tE/F+6DqsxsjgdvCvW1XZ8UQSAA4oebEBw5j8clH9EvbMN8tpmfP8IRtt60cL
NTxmY1UQl5ziBJ+SPESdFafBaPUE9LJ5jZ4IovFT0CXvngwOSrSJxcJ5YEmy+tsZHg9/MBBUYxpy
054edYm9MVsikIMMC8XFzIhx2LBUL85wK6IdUmK/7jghrtHkAGIqjozdg4HB0hKQh6cLPuKWpM/3
c2eZ+ecFj2yTjO2rl4u04IDxgTVXDEIj/Olc0RKQsaxUTpSL316L93pMcSrIBsPw+XukvhpM89BI
AgRGBA0loJ/JOV47WX5ziL5g7luq6j8QPv57K912wm/wNm9EzFEfpmbsJFLgm7FH1v807E0GPCSK
oQqrKqltg2BHBxTX31vphD7ADV+p5SvWGLf6zNhHqmvYd0J500lKNlgHTWgpUwH9mE0eqtsWGbzE
yAc+RSi7mP1OoWkI0VovGTI2y9euh/2CxOGLNJrA3iZrglvkMfA4UYpZtqrrP5Lcbx+ecoA7KxRU
pmEu5OLcoCVQHTpVFCZ5ScqnqV+UbE+qsEAY5GChBlWm+yUOfQMLgulGmkC1M9kSUAA7ayTFjHtK
FtQv1qFVE+AIm3B1e0GDI+SrrJismW+6/GkVjDyKiJagU+4Xyt70mBzGsm6027SjWXLruI8g+rzO
tMKa+VHH6VNc411opQQamDd/hN0qJWxz3jW+6PeUCCTRdh4huXuVhGNBDQZZlfsb9x/M23Hh3/8k
MNBvuyCV4VVew4Y2i8ivO9PNn4BhEeHm5drWFcg4ONdJW4+Rf5ktkOEMDrdJQMlWPoDW9kZ/pH50
f/Gr6noxMrVCwWeeVG/WMpnMNzEcuXybLA7CBRk8lcD6QYns7D8i5B48tN3zTV6+z5tJXytFQZlS
4VoxGF619RnjLjlYA74DHj5m0OL3DHXenPah2qoA3k7G8riGWVgNAEF/bpw/ybbHriVo6CoLtEfN
n5NsneMjFoEQE2wHdScxdC/L9xvwXbYKH09XYddP48D/tfB6zPSHpKiNf7xNAXhWpx8ScYhVND+X
jG7lI5XqYO1du7I3E8Eoqxef3zhD7FskG/yZJ4D7hz9QjeMFi01IccdL5iO/dwnGS7ElgJusw0ES
y7HhY/O/glyZvwJwQwslHs8j3JrkU1gdw77xSqPlib+Tr37cXWLJnLcD6sCdk3rTvcfY1TDQ0ksh
PkkQLKjWgUDlJmSbhlElnCENeaKcU1yGNqCH2r56FKFTXeWeByF4lbBW4kepNP7+2IFyDCoRc8d8
RNkEgAddI/YEhqSX7P+CJO/RuWZ3mw+VUcJq8gQ2sc9t4dY+mNksDBQi6NV9heJJJ5ahrTOiYrRs
iIsgTFCpiv9as/m3M/hbDpiBGpNgmeLEquSk+LGbgWD6ENyodkNTKPsHYtPnVerCMli/gmPA//xf
h19dR77YlNcj6rFDnfbepPFU8HfhF0Mus7qaeHiJbHX7JJ6pbvetDq7vKp6WLv4TnaAX0B7uACeq
qByAbneCnbSbT7HLlbVlttXCPPf+h6f6QjiIsE5WOvIHuAr7E6Ofqy3DkKFMnadMrU0AtTWRGjlo
nJTKVkhXvxkjEVSm9x+gneMhh3oCLVsbeWeXIhWWAqc59DLrRu13vcDID/ntrTonR2DywOwB8lhc
xiYIzivy8lC3WB4cgZF8CT3GDR5gATNCeGSXxHbnJq8MUcVzqfzlw0NNhb61q4FSDCUoO1/o8jlX
Y7PzJ0XpS0msWuYiH+Cwm2BGr6MqlTysFa1Xl4bcG8MrhtDFoebu4Oke+kMnH8+wjFIaYILxKaej
+H7YtnD7AYmIi04Tj6PB75iJNDmqw1srIUTIeho+4WVyWsKzdFnlrYW0SjtgGKLdQsVGwQU+odxR
yx0M6RfDzgcsHZESML/SakbZUfX+lyqMxiq0WErpAL5XKtCe/3RfM2mvAcj3Pt7mGlPxbQBJazu3
O+msa9uCCaRq4WOkduD0HVLyusABi+gHG3n3zcZ9MIOnz51p+aszfgeBs+OEwbsUj4xYCD6IaS8V
CjDHJgke5My+vI2ZkhVAVnYdZAQDXklJ6Kt7Yh2Ye5TMO7ZImdoAjfVhYqnpMoHDJQ/tF3VewhOI
suDQzHzWNUYts3KleO4cDUhdOIDZF6hwta7OhwZ5EojZmD/zkC2SQctiNOJDdu8LlL9JNWcSKYxE
tBA+ZfLdJujikqExiZK929ZcLkvjUNU+uLsdl2KhyItgdD/W0LBgfjCaLRdgz5khsidxxuGjlALu
HmZyvKr2cVL7ndsx7DvOzsmnb3IVyIosr1JS1X7s7JPRECUcU+InFHiEHgKpjAUXRGGPLNaXgiVI
iFXe4378UzT5kWGiS7my/HEVVQ6C7KIgJ5WBYPvq8KysCGewFSu3/Wp7lXDUPpTfK2UajdfJhbOl
7LFVN63QWBVRKMfLQB6eAsTI2+GaVrtBiMmMoT3/OKx280ZI5+Ap5SuzKpqwCivWzTn78VrQ50gj
WFfYeeFk4UoKvaxQ07hzxSeL5m9FuPyubpt6YVUdS6JfNQem7Qa/lVZ/GA+gxpv5Ab2N1m/UrW3f
6Wq/sC1bfCSlgOWj5BGeSCcLfh8G9Aq8MaByCbMH7GHM4Zigemj/ZoQ7moVBCnT1jTDA4NxO6cQl
iKiWr9GiX3LT+GHHczEp7yGtA9efLIpGgAjAdIA1zdm+CEd8aeJo55Ca6Up1UxOBHuiGI9YdH0ai
5bm1F5ihMqUCuERGW1oZKPnC8mQFC0iOfuvnL7gfFvYjn26hImKgzy3F4AHR3KgILE4MiTwqe2XW
aIwye2WiUb/NG26GXTEa4GIMheuAPrUD5gbj+13BG3wElczVf8Gq/7Jl96fZcexDf+bFSvqyGR3h
ZOlY7XX71i+BdX/0N6KbqvRE3hqvDLFBbKzRsd00u3stGRECvy2IkjIhWSdA1fBiq73qlv5JYdzQ
BSipniqCg/MrilRO9m/D671NkEcvkurzAX351n5A8zsTHH7ukyHdXbZn0/1QCj5BnEd9WDQ0yWix
ZGa0Pe7mlAbgBYQJxVqepvSDADniUHawSL4S3a4qve8qa6pkRRhItNcYAWjcqboNbvEMEDOIVIeu
KRKbbyjEKpEaiUPeTf7yfsumXN8vfy3dtPtTdG1cT0Q4dj9rQ6ZVVki2AYAixpBO9MgOrGCI7Uk6
6Vj5RPKQVoV0sdtHLrz7KTcbDEUL/71xiLGvms8rYcTspdLOufthTuKYbUDOe8KPiOWqkUhZJcbf
1Oz3dGFT41ciJqwcbSolx2MxFhvGESE/j18vRfcE2EI0qcuns3aApjxq0nYeW9bLtMJbVkfsBQQ7
B7/ru6WgODTVaaHlS8+IHvxw9WOfBYM0kSZWFBcVBJQZJD36ud+T5PmxcguIacslBTQrPUfXN3J4
CvCCUrt7jI5+5Io/PZhPgPH2MVreySkhUkBExaIa72ADuFqAdFOjsZPKIeKUukOACp4Sa/Md4UE8
iW8NfTfkaOxWuaX82MJ4GhztJzcVKzBoucGcQ13OMbMS6aQP0EmMnQjFBPuu4wfGd6saotGJXCZo
c7krXYtr8lUCUnhSBQJfwV7/ZOAMz9cfDLOfRqv3C6wM4/gd0s0wSw0AiKSwR5M030WSqeoAdsZV
1HvNb5emu0Weckur/iLT6kZrZ8lZxHCvT5Hzw7VKCes11qvSxaUA+ZXB7YVZSH1+390xqWKIZKYv
TUa2wIfLSLBM5OJ6TiUTwG8jlrBZiwbEGNn3kObd/ZEAWqFPVynQFLmqPdLkWQwoXK8Lf2T9oQLU
PpRL/0YQ7EexN2tRytDkJTwXV0TfISzvKDQjkHY71bdu/jb82Cgwk+zY/BCreNpIrCHIwjOGRhrE
g3vkg1fCjGBU13/KC7U8TXxOjTKhcONZPkkuXR6k/nmHuItnvWFYrawkTUuqa7sXbjkcYRVpfjaP
vqVH8X6o6Hu4dMx0TXquLJQryzQgxY6B06NJuUP3GYBGfB7Sw+JjfN7EIckhj15qWqF/g72ubbLd
L4ZFU8PvaDmob6b+Wv8u6xa8vG2IZbSzCuwnC0tHvgJl1XmcuhRGQCPId0QEDI9TJvVNtK+YgcwM
No6Fd9c0NiIq7UENPSwQFqQqtO4wkwsxp5loSRWQ81ZTfgaPv07gkNHjwRo6fozV0QRebsOCB6fy
BFF/G1pt/1enYDoKLin8SEoILRI8IRVqzhM1sLjESNeoifFwuoLSKdqHkg10JITc2LQoh/CbTT/f
8PddCx+1o31S1PrP6W71JFiMu3csaNvWs46/D5J6a4eg5zLT8cRso3gGBm6cQbljfbp7mTp+yUoS
IbDlIbiJ9QjeEqc0sKF0IycFn+EjEvK8Me4Q9yqTClP/PH0XYdt+VfItC2/1w/gDJuxxau4q9Kp0
lwJr/Ov7ZfeYkzFVjZaeOOLTYz4wH2AG0SHGWjoP6xe04lFSFbSd5zFl8GILL130GfzX4KY83KPz
9MXxlDwM0BZsuZnMFOK3GKM7GamZSAzeEf3Y7nc69XuV4Ev2G/G3xkYZVHmXhtT3dIqOVy2++Zja
ydDMhyxOHaiBD/MU4KkMb4ExpLMfrav0R5K+ho1qX6NYm0/86Y2XqCwQfZJBqSBcFGxKCSe8JmcZ
fQngV1n/HCX9eKtINrJ+YmFu8MUWk0u1hsMNnEwSVZdOQB+VL+KtMoyaNtM/ciM/756ukBBROu9m
edmfnUvG+Yef20wZc5aWEb/vTtzrdmQYtDOC45ve5u5aFZEhIdaLkMnF7ZjFoSbSYGM6IcaV7oeS
mkP23j+skN5GH1qwcWyYQ1pZ4++Q+I2TNtPaslBt0wD5HlvJgSh+ooV7qoaCNWg1z4qu7exp48h1
4tJG2QuSfA5aj8kJ4JmJANttXLsGcEXT2XYzhcuywdeCk5pIibMmZ/ePVNOTtK5i4IvW09MhZaCs
bpW10ykITw3Cynw/dsbiV9bYXaMKoAXvUYuvCPo4WQ20frL2ESLza2l+rwambwg3MsO/CaGS0kTO
ale00Eelma4khdMwwcOLpeL+FrAvdXB5+xt40YofA6ew9BvBHQAPzgFa89QxLJDlVvSYgoM6jYq8
ChQO5rSDFlETQ6Na7V4QiZfYsCS8/dQDXsfstttTeGxeBl7wc/tPr9bmvjRMlmCIxGvQMxxcHqMQ
iFUNLuE4juDH9yceNdW0yzq6+ohTySB7s11A5He6MjTFXs7mMO0Eozmr54jmtck4aQhJhg/t6TIr
JeCyJGI7GPt9FjmIni2i0mM0yrC4Oq/5HI7SnRU/BUT5xv7LrFspKQPhlL5SuIvguuidAYerXPQJ
Sb9zGbo3CSfQ4HWyEYSXt1BbXdVlcbD6y/5h/d6TX6UcUUQxX8WreEYIk/fA85w6VvLBAkKSs4Tu
fV8hX6kks1z5QdX4lruBeaxU1+DjMeuBZUTYtJih7FhqCsDwB6RxuZlGS7Jr4FYCoISDaS9zD61g
5FFGFY4FPKk9HO9pBjbyaGtKlYxe/q+I5o6s7BJbLIwySPpwCzW9RGiVffIzEXYkoIevfla8xjmv
Z1Yw4kkbvH03fQo7TSLoAQ1IJV8GO1AppC46X8XAkNhmJEg9CGtXq4c5v1B37xseP7uq/08Pe5b3
xHX1jKr1+mw4iqONTZLcgTlvbwULl35xE6BVtZFX0urrg4GVc8hKDgNphBG07+mvwYI62gadw/A6
vCuv0VBR9gylm2jexNt2T7Bajq254cDxFlwjaDImvmweCz1IXjN372zjrFetEZHu/uCAn8b1o+i/
GUeE9PQh+RWOhCDdzmhUE4hfCGwdyeb9b+VuD6rd4JPlOZwldeUVZjS9npwJrLVG9RU+yAzyGywB
H60z0GsghJLG6XTFkaOnrIQbWAwqALI5hJIaZQckCnBFrNTWPZBIwBuZF+E3voblzU9MXxf2Jd/M
jWzbaqZdskpSgvj7+4mq+DtqtSqzSVdGXJcVOWHgFF3dUQH0eP6uJTZaeyppP0TWdB9+NhsizfGH
+w26Q/hnSYchwMQhhdstFU12yiMmDIcZbaY+pDckzO4VjfIIxgIXzVzYOAiTNdP8gFP81ZUtqgNi
MFyq/vq1sZf0VuuniwD5xoE9TB9IjCLaA36D3/QVEcKMwJ+OUaYh2wQmmfBkBp57O8XM4Lz3KadI
dJyC0d7dtfwv7EOpT5OmF/XsfB6rlpSD7oeL+bgKahiuMOkow1JwafHtObH+tfWOYOUioOsLi/sU
lHnjXPLkIyWLl3EQ+S+sRZBvlmv3PMx6MNl4bMUG0zVINPKN6R9u3B5H8Pzvpfz/AmPONG9U61O0
GdPUWOp5FcH2ePadVK05oL1+/7gFQQozE0kBtzPAybTUG9NP6zHDMlXBaCooHib6Y9GYBNishfvm
GI8dL4mUoFBhwBLEPI65W1Xsy4ugFAvub6TILPVXkbwzpOvh1VxksaE6avG4TtzgLqz5Uuf0yaWl
iCOu3Ozy4Ik1YIHmM3+KhhO3Nm+JYFcNgatJX8ywbqypcmOplZXzpWiL7vMJ9+seeCt0pYKkJVMi
1AxbiMjcYrB+kOMX5TgvkrF5bPVz1zmgMBNjeVgNCW2YsojmyC/5aloc5HjGDORSFP0WM8S0xyHO
kIVu65WZlPUQbwjJ6dsWXYzjr1jeV25lR9WvTtW2vp/MEQIgjMmWyEdmQX6Pzzm1qbzeuRYjZT0l
5dHPSJUxz0FQ2+IX6CneB8fQaLhADpT23LaVdA8o2aFKjlsWdGRzUsP5Zqo0CQOqhhrLEb2RsAmH
PP+VhKYLMnSt3aAOUEebKKWRlKsbmopBcE3UgHkP/I0Wrn7RkrRqzUAEPM6JwKLwVr3i6ecUGMVz
7kXgyTsiiKzWrAiEHwXtsbCwY4NnQ6VkmZpIsLyqMZ5FXxdpvMJq6gBznywnsrMXpKiOCbd0b2Qm
6BlPssXSbfnegoFHRWred5d7PWswn2mJ7/Lyd3W/gXfIAh2Yv4FQ4fRkWVPEFaGeHn0FmIN+S8Pv
5bQr2NPK3cbOXezcQlBJOw2Nr7fkNdJVqSxWVqgf+Ay74GJqH9Abf3euZOx/BKmmpc9elKsD8FeH
mdTSfllB/DoDT+gxCfepHcpG8ZA5vtt1U0Si0VzQP80T60oOE3FhAd91GriI3iQzEng2uzwsejfu
GOR4ylipqWTbutgnqaUUGp5Oxan18E61FEmfvetBbeK86Cw4+2aDuFj2Lm74jkM9KxqWZk2acW23
rIyYeupF7ddkuwIpNYCv2s7JNmZodHU2XuV0p+m7nNHOaxBrEhtWltDiVnwUhqz73h2cA5VEakqQ
uHGcSEf+qjinIBkJdINqxEs8vxcN2eB0mY0JDTIYHQzqNWvGeSwrRFN/nS2od8/JhGTQxfz/gIj9
SYSTswPKotVXt0V+ZJFfZU0rn0opNyQuuJfxaOqHkKtGh8T2doDCGUedfT5MkmhGA+xTjv0EXw1t
I346opCTw1+UmRWACRTBplO/xR6OkmUr3ywm7lViMbZjkl4a8oAPB0ZqsQuSci7IkQUkjY6OZ/MH
0CqD4WPOFlF4vqlgfYegVh9OdbX5wI258QF1TvH40YYPe55BBZDE8V6gupriyDDrcfwPINWN0hEA
CN9sfqi/icaX3wK2AWfPMTYRBaodlkXiMSTYZdTDXpciZZzFfxIwWxpl12t2OIaKdyTOnySvhyoS
Y+6ZNIbQ4TjPPIVI1Z8yHK7/3zbmVkxeZQ10GISV7hrolTHAfcBaD7zUP/K0JbR/iX6q2kHcA5ar
pbXpyHstU78FsQZANcbd5ExfMUnTofXbhiJJcXZBu82RXj7bn4B15Q+9oCmhA0XoBem2En1kGdAY
24EDHlmIBgbW7h8CR2VXA5kOhPkD4NTs0W8uI7us3SGG8JPgkeVp4jmCYUIxQOMw8b81vXmhfEqV
U0cGt4nMSAP59np9Bdk92dD80WlceDdnWOTaZLa83oTyLHaz43/3ZuPqh3Xadz/fpJeHx/6Xt6Rh
uYnGvjN7YxoC8D7QT4xztNeB0dFP9jzfV7C4XwTjPYDfPeZhg+KLddxrqZdEt7KEde8QGwXxr85h
FkGGMVzJ3ljgSFFN9ab1D4BPTje9VrnNDm1awwwF/sNFl8NcF75D9gLFCQlsG/AsRqyj/+fGwjpp
mvyFOUsHcowxPYcVRkYnttLiylK1EWs0IPX22wEIdpTjbmSSPNGjG5/GuQB1vNINg1wIRkVnqfdO
t6GYl801wU/TGXwLL3XuUe/EEgz/0a1dJo8WrRJxKYk/nnLuBH176wkeaLh5VEUoDNc2sAXE0hTm
7ESyr0/uJBJX0bkWw7wfP40azrAKmRdVm8j0UYljAV9flDOgIDwh9jRjo5rcEyRYwwm2lHk2CLAV
j/uVtpiCf8XOuEkXeRB1AwWCFv3X/piohv52Awvy/XHpazBJstqrfw9gWrna8TkRc2hZ1i8JEb/U
qGAhVJUvwxX4NPNnrH0IpzdOfcxFn5XxOZDopjlUQLJX/DYNFeOGSs8bfyYIj9dPMkoMbECNDiAJ
FKQBGcNe1TXDTt79+LWYP3+CAYe7U7MFTSDOhATe95RIy0c/zUlGnVyTzBJFw3yQinLXmfQMcntw
A6ffwS1QOEfVdvAHqUnFZNSg7M6BqH/ytisKcAc9+8eWAPHXV3EG+JAYGo0JIzBwpJPAzsotxbI4
p6GwohakAV/2oWtFnHM1b0AA+lUjcwc/WSDnIczNObXW6i6s4b/2mijdVg03bgB1kEYmZZKLDZ7g
kiV73cjYmOR3nNABLZs+I79v18f3VCdDOEzUprd3qdPpJgWRMAHJI+riIAmbbsO+DQ3oX6t9Ysom
zo5cCBv4xQ6m3xx2dUXN0PupHhbnpKquitlqgrr6C1mEXPu1l3+9zPF8TP1NdGYBEqBZ+loHf1iy
F2UjRSegiUtzrPglW3hmrVkiA4iTMZ34iacTH+YyUMfA2/REluaJjIFDx+lzxcD1+eI4MRES2RCr
k24Ohl+mG+rn+7IXe73gqPQwlyvBY6Q306sSeRegfQZhCvjKjTPd+xYZfvYPdXtMTi8vYugc62Oa
oYsfRLsKlWGp/JguoLal3umf9O89Y1o88MDn36rYXxu6lvDOC1JrV/rfyNo2zasXRy/qJ5waqFgE
H/CY3v/jGPyDq/4tmM3pBZmWwS5BHYyV8VMh+Yb5fI1m1TBrzk1tDtk4jlA0j9/1xxGfCPL245sa
22ydLlxdwEhHvv5m2xXXUCEE4AwxD3zWbBvB4eDRZRDrwC1Rr4Bk5B+Y7qop64MkKp6FjJd/UEwW
sOPx0vteYC+bfOKmQZ/sjYAgcDY1CGR6axRienrwsW7V4KIlYRBw/csGFPUdfv80TW/8C6jOngVg
VymhR7jMzN0/HuDgTBV9osaomia0ONlaOkCD3NoLjDVvmplqOAcn3SvMNL8G6hKq09FU4ol/jkoR
9RPfOtpY8nz5i6aUt0BBhyd0SGNIS0oqX9XbC6OjynrWrMkvEkc44vStU2SMBkls88oFEWTrzzbt
L0EmgU5/PLhKyqDT0EYqcppTxLP34Og/78btf9a30Zm1GWmT9c8Cv7wVqcCldJcT2dffrBmnsV5l
1EAqRIKwFrtbj38lt+o5TuFMpxd87bLhD1udYqAWEck3UgUeoUbmbUY65wiQl3S/bDegXUASpMEO
v7T2MZITuUDXG1Dr3ySvB826Opo1ywsEy2TI1e2crSoEe+CZVIZZ9NXWyl7OPsanyd2MIn6fDgoL
Wa9oi0ht0bEk2WkZ0H6tzspofAZH5EJTOZMFm2pux8m39Dp3xJ+fJxFKI9B86VLpiW5bwWDRoG/W
HT7MjzxFQ8A0MlmCZuz+mdkY96x3MH1QuNIeYPIRf4M58uP96KJm/w8OiWHZQxcxzx18w054Macr
cU72xxHecFYjOZAp9ox9uLJpJuQwyOrW4HQSNOnqfAFH4LRwLBytMi0yxRW1sVxmnCwLtmEg0kxn
bfusKqM0KiBgA/fmAT0M91gK2Kbqk1PMExQxyg0sBYJxfCxoR1Qpu/cvYz+6pRQhLbEdTEFvZoBd
/CX+XAZWiAe5TpxnkAjC+fzzoQAkaSfQhRpqttCQa5A1nPUr7c6vagWtT+eSkROMP61ImW7rG/sp
3OoTgMHDzAea2GykmnxVeb5o6d7UUKElnD1qwA3vafXtr2lTE8p2iu4lBx34rof09tLar8yNIkAq
SmNXoVAGTeA7o9Tbwl6DqfYD0G+lzWGYohzot59mwZIdKwUEIODZlubVo/jbySTXVKoNO9PLMEva
9z1rHTKv2D2miBa5mUCQlUT/vrzwIRSv1GEvuaCwr7I1/xGSv0G7u+rkxocWmbj5nJZqZ38Nlobo
DoVB3jhdqT2u0QpgXFzEVr2g/aSNkvGh0Y7Qmq6SlQRvqKqC0MgI3ZIxWzkQISp0eoJERxsw1Dae
X5hMEsi/rv5zpdnPuC5ZV7dgUvE1oAkskkaik+ZTzp7jFzez4EwZ1J0ztIYv3nERRqH7SxRtK9OV
C9ouMhrF9JwBu7h6UZ/NTh/43wTj9VwjPmJDlI58YnCAjbzbYkPkpo0zt1pzlEKz0v9itKNjYVCb
zaKsE9wSNVaaj/9bjsyj7gWG9J1Ib2ijfwu8A3WHPtZBkl82cMb3X9NFLyf5f0ITirJjuJ3BYldX
zp1DW9BTMtU5TukcjbOOPdcRa11nkpCPdGKyKssvHqqB07aic/9ctjMl0g/lYoiKfSBpr//rpQRz
MxC91NBSU2PgalluK7uq6hYHmUZTj8wvUR6zgUCj0JOD4HbQyHcH3P8AhSrOUqOuVhx+EWYDlkjr
QIJk4Eale7sLsMRbYJYZQBLgxSaC+GjF2bZUoKpUyZyn4w3Ofrjox9gMGK7t8u0JZzfWoANWGczr
ha6tL1xGALcpXq2aruHPcn1MWuRyaoA2OfRWvMbUXLCE0i8262LfiHtEliYmRVdFpR/JDwKhry+U
OxNxoHWM8vPOu33XHgcllzCEeIdgNv7AswnQI0rFOW5iEp1Tan31nQNPtgdveCebUeKUj+X9x9Io
x0JqsQrkKDfSDDcuNZ8L0Oggo7Jq3eCPn4gTYDX6Ux1Rdk2AGNWRnocMtetilZ8Vg+xP705YkYOq
+wXty8BMuZf8KaNK0G7FEc2A+PPm8nr/Yhdx0/lmIHy4N5YE8E3Vd1EHUFymPO3YB0jrbbEwOR4Q
aT1Y9QhwyfdQSQpR+KG2NzwPHjFmttcPxMVyR3Unm7ppVmf4+KRkPZ9Ns29LmzSGOXmxE93Fwiw7
gk44OOZ+hbR6+jdY8ztNOn8YntrxHBsvVn58AYxCve8QqKTmQqpJQBYH2XHllEjNNhvHXUIJ1qp5
hfp0TJ450TOTwb+PZFl+ARam5Ffg6Kyp3U007gXn5Xkb7PThltNsfj0H9sfVvSNmfu7MNjVkzahw
riloL+6se2EaB029sx3uKZmCxGTV5SS14yPu1FnDPuq731q0F8WVRM3VqfG6gNu9RWTkkh0jIrJ8
AtTdQ1YzdJ9lDThq2jVBNI2yWsIT2E+19ON7eOLV+QJ91DCKZqbpC6MNp9dnTyiZze7QEtT/rvfY
+Z/g+CvXifOGRlYc7jDLx2yCntY+hZuQ5BMqzx4mKRKLNEmK7IThOtyDzcJ5/16PrD1SvGh2KSz4
5xcM6+rOcjUfLNdYGtLtHeh/kei1Mcy2mwXKeap/IUSSl+8VT3tX1LtxP12nfr0dzOT2uSrA2wa3
/HEeWReWV+Zj36LlYrenz8hXfYjzMs2vRpe2k2HAi9ymYI+pVEWXmR7dLJcQcXT0Wt/GvFvNgjYT
peWGe9+Ds/W9c9ltxqHJEvjEAofud64DUDXe5xLWkdgnJBi3+SnsGQdIl5gwwfwYoUKzj44lZIu9
JKgG/eWwztyd9rUGoMofDZMpMgEoe97q/xj1pZFRrz2WJtOmVp+aPpnVJoblsGenpEmHSirTnvVs
mVyADsTRYKi9T2j6UsXa55lf5+Nai0Zhk0Cq5ER5RXPcHBnFUdRmLdmWa18Ij+8QJEEnr0F62Zmw
7PXIuKFzAdMnhO8JsGLYUKhmcj1w7m4ALxULWMvtlFRUCOA/7dIna4/mcAuXXbP5J9BKfWC7CqD8
uWdZ7t8CNVbHOGaumQPgquc5Y4aN5kjtksJA5dPIDx2kFGa5uyBgUfSYTwyq0Ioy/NtboMKk650z
q13iA+0o7qWQPaLyzu9BOor0NIvfPLv6KwJ6AE28q/iWf/VQr32wxYg0vtZyRH+1cxtAUp5ZT4P7
H6hXXgvkO1Sx4ycssh9fM5AqnSJEBOBVkU297tFPsvpNcu0mxGVEPEQmU9pNFB+V3bXwm74eXN/w
UcM3dvPxsF5foe2RbMX7UEBthpTnZV/zKvFZakEBzZ73WTsytu4okHqLsTJij6n9PfbpPYxMwDY1
g5764vGg8ocXcrX8/yjQOD6HPXhVy5CBt44zjDZF9GiwEWaZvs9xGKeZkEp46Hk4enQXMtYhiMmw
l1NasRAdCswGNGIbgsi4K/b0ZKNmDQDpRAgj4PY7OLF7tJJw7PTcOazBL2EklLkX5+doDIqjDVMo
7BK9gkMKqOUxT7/RGvdczRY5kZunSHypUDIsitbK0rcSHsd5XiGe3VQQ7ljDC7CITwSLGBeRMPGe
GfBVCfGsM0SpdMXxqnKv27KOXK6rUnb01Nh2Dsw8AHZUbbmU+tZK7UTMainm2TOi7AOlrTPFRYN/
q/+5hd4rQpFVKIj2+gZzdEAIbmqVTaEuWBcS9AGWUSaGZ/PVl7cXL4Nh1mBMS4h2JH8qpykB7hcU
3Q4bkajm5vOEU24yldLD/+8WfnI1gST1dnqQcen9gq2ocAorH2hkxY+DK8M82LMO+CEf9ieqbDea
14gnc448t1X9kB5RFi8KtwOgw86P5P8uiZ/1IOAxXJZ65p+NbCiIrl1xDeRNvkjJdOp8Y55zud9Q
4al9T06F+1RqcjXrNc73TN75bLdeCpi1lmdDBWwZKssh0PEYJ9vTmUSTNJ5Y91oHMWgJAyEi9jg1
ieypCQV04bj2yAyl+wkU1YMJsTVyxpyCvmxOLEDi52TqKthKjQo+E7pfJIxel9A++Paeg3rDCud0
9iUGldMjoaXXNXhxIA8w+L1eJxRyxWV3F3dNVJUjXP61IREy174EkxBV14/eiHawIPGKySf+KjPq
pTwtlpge1pDcnLWHVJAIP5lp1VOdlqkOAvo9TY6sx7sAeWTDLgNdcC883x4XtlJ5G1QuhpiuVfKw
negRoaQ2eVxUh9pSV+6UoYxtXQvGDb9rpeIjLLfwQ/PEHcI5AwJwf30ojfUoz571Bq98Z/NiEPYO
ZBERWIFl1tcj
`protect end_protected
